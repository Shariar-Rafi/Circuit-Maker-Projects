CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
216 93 1364 691
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
426 213 567 334
42991634 0
0
6 Title:
5 Name:
0
0
0
30
5 SCOPE
12 685 592 0 1 11
0 7
0
0 0 57568 0
3 TP2
-11 -4 10 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5130 0 0
2
44824.4 29
0
5 SCOPE
12 685 478 0 1 11
0 8
0
0 0 57568 0
3 TP3
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
391 0 0
2
44824.4 28
0
6 74112~
219 265 327 0 7 32
0 7 19 2 19 8 48 12
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U7B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 7 0
1 U
3124 0 0
2
44824.4 27
0
7 Pulser~
4 61 341 0 10 12
0 2 46 2 47 0 0 10 10 1
7
0
0 0 4640 0
0
3 V13
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3421 0 0
2
44824.4 26
0
14 Logic Display~
6 346 123 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
44824.4 25
0
14 Logic Display~
6 636 124 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
44824.4 24
0
6 74112~
219 554 315 0 7 32
0 7 18 13 18 8 45 11
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U8A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 8 0
1 U
8901 0 0
2
44824.4 23
0
6 74112~
219 843 302 0 7 32
0 7 17 14 17 8 44 10
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U8B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 8 0
1 U
7361 0 0
2
44824.4 22
0
14 Logic Display~
6 915 123 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
44824.4 21
0
6 74112~
219 1131 291 0 7 32
0 7 16 15 16 8 43 9
0
0 0 4704 0
5 74112
4 -60 39 -52
4 U10A
19 -61 47 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 9 0
1 U
972 0 0
2
44824.4 20
0
14 Logic Display~
6 1203 121 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
44824.4 19
0
9 2-In XOR~
219 400 297 0 3 22
0 12 6 13
0
0 0 608 0
5 74F86
-18 -24 17 -16
4 U11A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
9998 0 0
2
44824.4 18
0
9 2-In XOR~
219 693 293 0 3 22
0 11 6 14
0
0 0 608 0
5 74F86
-18 -24 17 -16
4 U11B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
3536 0 0
2
44824.4 17
0
9 2-In XOR~
219 1003 280 0 3 22
0 10 6 15
0
0 0 608 0
5 74F86
-18 -24 17 -16
4 U11C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
4597 0 0
2
44824.4 16
0
12 Hex Display~
7 1284 271 0 18 19
10 12 11 10 9 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3835 0 0
2
44824.4 15
0
5 SCOPE
12 165 322 0 1 11
0 2
0
0 0 57568 0
3 TP4
-11 -4 10 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3670 0 0
2
44824.4 14
0
5 SCOPE
12 326 279 0 1 11
0 12
0
0 0 57568 0
3 TP5
-11 -4 10 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5616 0 0
2
44824.4 13
0
5 SCOPE
12 614 268 0 1 11
0 11
0
0 0 57568 0
3 TP6
-11 -4 10 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9323 0 0
2
44824.4 12
0
5 SCOPE
12 893 256 0 1 11
0 10
0
0 0 57568 0
3 TP7
-11 -4 10 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
317 0 0
2
44824.4 11
0
5 SCOPE
12 1184 244 0 1 11
0 9
0
0 0 57568 0
3 TP8
-11 -4 10 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3108 0 0
2
44824.4 10
0
5 4023~
219 533 502 0 4 22
0 11 9 5 8
0
0 0 608 0
4 4023
-14 -28 14 -20
4 U12A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 11 0
1 U
4299 0 0
2
44824.4 9
0
9 Inverter~
13 428 528 0 2 22
0 6 5
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
9672 0 0
2
44824.4 8
0
9 Inverter~
13 426 582 0 2 22
0 9 4
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
7876 0 0
2
44824.4 7
0
9 Inverter~
13 420 621 0 2 22
0 11 3
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
6369 0 0
2
44824.4 6
0
5 4023~
219 491 604 0 4 22
0 4 3 6 7
0
0 0 608 0
4 4023
-14 -28 14 -20
4 U12B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 2 11 0
1 U
9172 0 0
2
44824.4 5
0
13 Logic Switch~
5 152 244 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7100 0 0
2
44824.4 4
0
13 Logic Switch~
5 441 232 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3820 0 0
2
44824.4 3
0
13 Logic Switch~
5 730 219 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7678 0 0
2
44824.4 2
0
13 Logic Switch~
5 1018 208 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
961 0 0
2
44824.4 1
0
13 Logic Switch~
5 144 399 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3178 0 0
2
44824.4 0
0
51
1 0 2 0 0 16 0 16 0 0 3 2
165 334
165 332
1 0 2 0 0 16 0 4 0 0 3 5
37 332
27 332
27 318
123 318
123 332
3 3 2 0 0 16 0 4 3 0 0 4
85 332
227 332
227 300
235 300
2 2 3 0 0 16 0 24 25 0 0 3
441 621
441 604
467 604
2 1 4 0 0 16 0 23 25 0 0 4
447 582
445 582
445 595
467 595
2 3 5 0 0 16 0 22 21 0 0 4
449 528
507 528
507 511
509 511
0 1 6 0 0 16 0 0 22 33 0 3
267 399
267 528
413 528
1 0 7 0 0 16 0 1 0 0 23 2
685 604
685 604
1 0 8 0 0 16 0 2 0 0 28 4
685 490
685 517
684 517
684 515
1 0 9 0 0 16 0 20 0 0 40 2
1184 256
1184 255
1 0 10 0 0 16 0 19 0 0 43 2
893 268
893 266
1 0 11 0 0 16 0 18 0 0 46 2
614 280
614 279
1 0 12 0 0 16 0 17 0 0 49 2
326 291
326 291
0 1 9 0 0 16 0 0 23 29 0 5
328 502
328 566
394 566
394 582
411 582
0 1 11 0 0 16 0 0 24 30 0 4
402 455
341 455
341 621
405 621
0 1 12 0 0 16 0 0 15 49 0 4
345 164
1340 164
1340 295
1293 295
0 2 11 0 0 16 0 0 15 46 0 5
636 172
1316 172
1316 313
1287 313
1287 295
0 3 10 0 0 16 0 0 15 43 0 6
915 157
915 153
1308 153
1308 328
1281 328
1281 295
4 0 9 0 0 16 0 15 0 0 40 6
1275 295
1265 295
1265 352
1328 352
1328 140
1203 140
0 1 7 0 0 16 0 0 3 21 0 3
554 179
265 179
265 264
0 1 7 0 0 16 0 0 7 22 0 3
843 179
554 179
554 252
0 1 7 0 0 16 0 0 8 23 0 4
1131 178
1131 179
843 179
843 239
4 1 7 0 0 16 0 25 10 0 0 5
518 604
1253 604
1253 178
1131 178
1131 228
0 3 6 0 0 16 0 0 25 33 0 4
213 399
213 639
467 639
467 613
0 5 8 0 0 16 0 0 3 26 0 3
569 340
265 340
265 339
0 5 8 0 0 16 0 0 7 27 0 4
844 339
844 340
554 340
554 327
0 5 8 0 0 16 0 0 8 28 0 3
1131 339
843 339
843 314
4 5 8 0 0 16 0 21 10 0 0 4
560 502
560 515
1131 515
1131 303
2 0 9 0 0 16 0 21 0 0 40 5
509 502
298 502
298 412
1199 412
1199 255
1 0 11 0 0 16 0 21 0 0 46 5
509 493
402 493
402 423
603 423
603 279
0 2 6 0 0 16 0 0 14 32 0 4
659 399
982 399
982 289
987 289
0 2 6 0 0 16 0 0 13 33 0 4
362 399
661 399
661 302
677 302
1 2 6 0 0 16 0 30 12 0 0 4
156 399
364 399
364 306
384 306
3 3 13 0 0 16 0 12 7 0 0 4
433 297
474 297
474 288
524 288
3 3 14 0 0 16 0 13 8 0 0 4
726 293
808 293
808 275
813 275
3 3 15 0 0 16 0 14 10 0 0 3
1036 280
1101 280
1101 264
1 1 10 0 0 16 0 9 14 0 0 4
915 141
971 141
971 271
987 271
1 1 11 0 0 16 0 6 13 0 0 3
636 142
677 142
677 284
1 1 12 0 0 16 0 5 12 0 0 3
346 141
384 141
384 288
1 7 9 0 0 16 0 11 10 0 0 3
1203 139
1203 255
1155 255
0 4 16 0 0 16 0 0 10 42 0 3
1070 208
1070 273
1107 273
1 2 16 0 0 16 0 29 10 0 0 4
1030 208
1092 208
1092 255
1107 255
1 7 10 0 0 16 0 9 8 0 0 3
915 141
915 266
867 266
0 4 17 0 0 16 0 0 8 45 0 3
782 219
782 284
819 284
1 2 17 0 0 16 0 28 8 0 0 4
742 219
804 219
804 266
819 266
1 7 11 0 0 16 0 6 7 0 0 3
636 142
636 279
578 279
0 4 18 0 0 16 0 0 7 48 0 3
493 232
493 297
530 297
1 2 18 0 0 16 0 27 7 0 0 4
453 232
515 232
515 279
530 279
1 7 12 0 0 16 0 5 3 0 0 5
346 141
346 164
345 164
345 291
289 291
0 4 19 0 0 16 0 0 3 51 0 3
204 244
204 309
241 309
1 2 19 0 0 16 0 26 3 0 0 4
164 244
226 244
226 291
241 291
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
651 31 716 55
662 40 704 56
7 Counter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
478 30 633 54
489 39 621 55
22 MOD 10 Asynchronous Up
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1206 78 1254 101
1219 88 1240 103
3 MSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
287 81 335 104
300 91 321 106
3 LSB
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
