CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
34
13 Logic Switch~
5 128 820 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90043e-315 5.26354e-315
0
13 Logic Switch~
5 127 772 0 1 11
0 11
0
0 0 21360 0
2 0V
-8 -16 6 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.90043e-315 0
0
13 Logic Switch~
5 115 542 0 1 11
0 17
0
0 0 21360 0
2 0V
-8 -16 6 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90043e-315 5.36716e-315
0
13 Logic Switch~
5 116 590 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.90043e-315 5.3568e-315
0
13 Logic Switch~
5 103 312 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-8 -16 6 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
44796 0
0
13 Logic Switch~
5 104 360 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
44796 1
0
13 Logic Switch~
5 101 184 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
44796 2
0
13 Logic Switch~
5 100 132 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
44796 3
0
13 Logic Switch~
5 99 84 0 1 11
0 30
0
0 0 21360 0
2 0V
-8 -16 6 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
44796 4
0
14 Logic Display~
6 725 299 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.90043e-315 0
0
14 Logic Display~
6 699 253 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.90043e-315 0
0
14 Logic Display~
6 675 208 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.90043e-315 0
0
9 2-In AND~
219 408 905 0 3 22
0 6 7 9
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3536 0 0
2
5.90043e-315 5.36716e-315
0
8 2-In OR~
219 521 930 0 3 22
0 9 8 2
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
4597 0 0
2
5.90043e-315 5.3568e-315
0
9 2-In AND~
219 232 947 0 3 22
0 11 10 8
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3835 0 0
2
5.90043e-315 5.34643e-315
0
9 2-In XOR~
219 424 792 0 3 22
0 7 6 3
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U4D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3670 0 0
2
5.90043e-315 5.32571e-315
0
9 2-In XOR~
219 231 790 0 3 22
0 11 10 7
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U4C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
5616 0 0
2
5.90043e-315 5.30499e-315
0
9 2-In XOR~
219 219 560 0 3 22
0 17 16 13
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9323 0 0
2
5.90043e-315 5.34643e-315
0
9 2-In XOR~
219 412 562 0 3 22
0 13 12 4
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U4B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
317 0 0
2
5.90043e-315 5.32571e-315
0
9 2-In AND~
219 220 717 0 3 22
0 17 16 14
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3108 0 0
2
5.90043e-315 5.30499e-315
0
8 2-In OR~
219 509 700 0 3 22
0 15 14 6
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
4299 0 0
2
5.90043e-315 5.26354e-315
0
9 2-In AND~
219 396 675 0 3 22
0 12 13 15
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9672 0 0
2
5.90043e-315 0
0
9 2-In XOR~
219 207 330 0 3 22
0 24 23 19
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
7876 0 0
2
44796 5
0
9 2-In XOR~
219 400 332 0 3 22
0 19 18 5
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6369 0 0
2
44796 6
0
9 2-In AND~
219 208 487 0 3 22
0 24 23 21
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
9172 0 0
2
44796 7
0
8 2-In OR~
219 497 470 0 3 22
0 22 21 12
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7100 0 0
2
44796 8
0
9 2-In AND~
219 384 445 0 3 22
0 18 19 22
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3820 0 0
2
44796 9
0
14 Logic Display~
6 652 158 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
44796 10
0
14 Logic Display~
6 637 97 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
44796 11
0
9 2-In AND~
219 361 228 0 3 22
0 28 27 26
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3178 0 0
2
44796 12
0
8 2-In OR~
219 493 242 0 3 22
0 26 25 18
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3409 0 0
2
44796 13
0
9 2-In AND~
219 204 259 0 3 22
0 30 29 25
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3951 0 0
2
44796 14
0
9 2-In XOR~
219 396 104 0 3 22
0 28 27 20
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
8885 0 0
2
44796 15
0
9 2-In XOR~
219 203 102 0 3 22
0 30 29 28
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3780 0 0
2
44796 16
0
45
3 1 2 0 0 8320 0 14 10 0 0 3
554 930
725 930
725 317
3 1 3 0 0 8320 0 16 11 0 0 3
457 792
699 792
699 271
3 1 4 0 0 8320 0 19 12 0 0 3
445 562
675 562
675 226
1 3 5 0 0 8320 0 28 24 0 0 3
652 176
652 332
433 332
0 1 6 0 0 4096 0 0 13 7 0 5
421 812
421 886
376 886
376 896
384 896
0 2 7 0 0 4096 0 0 13 12 0 3
290 790
290 914
384 914
3 2 6 0 0 12416 0 21 16 0 0 6
542 700
554 700
554 812
400 812
400 801
408 801
3 2 8 0 0 4224 0 15 14 0 0 4
253 947
489 947
489 939
508 939
3 1 9 0 0 4224 0 13 14 0 0 4
429 905
486 905
486 921
508 921
0 2 10 0 0 4224 0 0 15 13 0 3
163 820
163 956
208 956
0 1 11 0 0 4224 0 0 15 14 0 3
187 772
187 938
208 938
3 1 7 0 0 4224 0 17 16 0 0 4
264 790
400 790
400 783
408 783
1 2 10 0 0 0 0 1 17 0 0 4
140 820
207 820
207 799
215 799
1 1 11 0 0 0 0 2 17 0 0 4
139 772
207 772
207 781
215 781
0 1 12 0 0 4096 0 0 22 17 0 5
409 582
409 656
364 656
364 666
372 666
0 2 13 0 0 4096 0 0 22 22 0 3
278 560
278 684
372 684
3 2 12 0 0 12416 0 26 19 0 0 6
530 470
542 470
542 582
388 582
388 571
396 571
3 2 14 0 0 4224 0 20 21 0 0 4
241 717
477 717
477 709
496 709
3 1 15 0 0 4224 0 22 21 0 0 4
417 675
474 675
474 691
496 691
0 2 16 0 0 4224 0 0 20 23 0 3
151 590
151 726
196 726
0 1 17 0 0 4224 0 0 20 24 0 3
175 542
175 708
196 708
3 1 13 0 0 4224 0 18 19 0 0 4
252 560
388 560
388 553
396 553
1 2 16 0 0 0 0 4 18 0 0 4
128 590
195 590
195 569
203 569
1 1 17 0 0 0 0 3 18 0 0 4
127 542
195 542
195 551
203 551
0 1 18 0 0 4096 0 0 27 28 0 5
397 352
397 426
352 426
352 436
360 436
0 2 19 0 0 4096 0 0 27 33 0 3
266 330
266 454
360 454
3 1 20 0 0 8320 0 33 29 0 0 4
429 104
429 125
637 125
637 115
3 2 18 0 0 12416 0 31 24 0 0 6
526 242
530 242
530 352
376 352
376 341
384 341
3 2 21 0 0 4224 0 25 26 0 0 4
229 487
465 487
465 479
484 479
3 1 22 0 0 4224 0 27 26 0 0 4
405 445
462 445
462 461
484 461
0 2 23 0 0 4224 0 0 25 34 0 3
139 360
139 496
184 496
0 1 24 0 0 4224 0 0 25 35 0 3
163 312
163 478
184 478
3 1 19 0 0 4224 0 23 24 0 0 4
240 330
376 330
376 323
384 323
1 2 23 0 0 0 0 6 23 0 0 4
116 360
183 360
183 339
191 339
1 1 24 0 0 0 0 5 23 0 0 4
115 312
183 312
183 321
191 321
3 2 25 0 0 4224 0 32 31 0 0 4
225 259
461 259
461 251
480 251
3 1 26 0 0 4224 0 30 31 0 0 4
382 228
458 228
458 233
480 233
0 2 27 0 0 4096 0 0 30 42 0 3
304 184
304 237
337 237
1 0 28 0 0 8192 0 30 0 0 43 3
337 219
329 219
329 102
0 2 29 0 0 4224 0 0 32 44 0 3
135 132
135 268
180 268
0 1 30 0 0 4224 0 0 32 45 0 3
159 84
159 250
180 250
1 2 27 0 0 4224 0 7 33 0 0 4
113 184
372 184
372 113
380 113
3 1 28 0 0 4224 0 34 33 0 0 4
236 102
372 102
372 95
380 95
1 2 29 0 0 0 0 8 34 0 0 4
112 132
179 132
179 111
187 111
1 1 30 0 0 0 0 9 34 0 0 4
111 84
179 84
179 93
187 93
85
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
949 76 1002 100
959 84 991 100
4 Sum:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
1114 40 1247 64
1124 48 1236 64
14 ID  : 20201058
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 30
1114 0 1247 44
1124 8 1236 40
30 Name: Md.Monem 
Shariar Rafi
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
949 141 1002 165
959 149 991 165
4 0101
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
737 912 798 936
747 920 787 936
5 C out
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
343 329 380 353
353 337 369 353
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
359 299 396 323
369 307 385 323
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
421 303 454 327
429 311 445 327
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
523 445 548 469
531 452 539 468
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
469 476 494 500
477 484 485 500
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
466 442 491 466
474 450 482 466
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
220 462 257 486
230 470 246 486
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
164 493 201 517
174 501 190 517
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
164 454 201 478
174 462 190 478
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
339 451 376 475
349 459 365 475
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
334 418 359 442
342 426 350 442
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
405 422 434 446
415 430 423 446
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
174 345 211 369
184 353 200 369
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
232 305 257 329
240 313 248 329
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
170 291 195 315
178 298 186 314
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
465 249 490 273
473 257 481 273
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
516 218 541 242
524 226 532 242
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
464 211 489 235
472 219 480 235
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
375 207 400 231
383 215 391 231
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
325 234 350 258
333 242 341 258
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
327 196 352 220
335 204 343 220
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
165 227 190 251
173 235 181 251
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
221 235 250 259
231 243 239 259
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
163 263 192 287
173 271 181 287
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
370 117 399 141
380 125 388 141
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
366 72 391 96
374 80 382 96
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
432 99 461 123
442 107 450 123
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
159 50 184 74
167 58 175 74
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
230 80 259 104
240 88 248 104
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
171 115 200 139
181 123 189 139
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
636 469 673 493
646 477 662 493
2 C2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
586 330 623 354
596 338 612 354
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
534 239 571 263
544 247 560 263
2 C1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
509 91 546 115
519 99 535 115
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
41 169 94 193
51 177 83 193
4 C0=0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
355 559 392 583
365 567 381 583
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
371 529 408 553
381 537 397 553
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
433 533 466 557
441 541 457 557
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
535 675 560 699
543 682 551 698
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
481 706 506 730
489 714 497 730
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
478 672 503 696
486 680 494 696
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
232 692 269 716
242 700 258 716
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
176 723 213 747
186 731 202 747
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
176 684 213 708
186 692 202 708
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
351 681 388 705
361 689 377 705
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
346 648 371 672
354 656 362 672
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
417 652 446 676
427 660 435 676
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
186 575 223 599
196 583 212 599
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
244 535 269 559
252 543 260 559
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
182 521 207 545
190 528 198 544
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
194 751 219 775
202 758 210 774
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
256 765 281 789
264 773 272 789
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
198 805 235 829
208 813 224 829
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
429 882 458 906
439 890 447 906
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
358 878 383 902
366 886 374 902
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
363 911 400 935
373 919 389 935
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
188 914 225 938
198 922 214 938
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
188 953 225 977
198 961 214 977
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
244 922 281 946
254 930 270 946
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
490 902 515 926
498 910 506 926
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
493 936 518 960
501 944 509 960
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
547 905 572 929
555 912 563 928
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
445 763 478 787
453 771 469 787
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
383 759 420 783
393 767 409 783
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
367 789 404 813
377 797 393 813
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
564 695 601 719
574 703 590 719
2 C3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
555 928 592 952
565 936 581 952
2 C4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
557 562 594 586
567 570 583 586
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
567 788 604 812
577 796 593 812
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
246 3 363 27
256 11 352 27
12 4 Bit Adder:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
947 107 1000 131
957 115 989 131
4 0011
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
947 90 1000 114
957 98 989 114
4 0010
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
50 65 83 89
58 73 74 89
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
50 115 83 139
58 123 74 139
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
47 296 84 320
57 304 73 320
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
51 342 88 366
61 350 77 366
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
59 526 96 550
69 534 85 550
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
63 572 100 596
73 580 89 596
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
71 756 108 780
81 764 97 780
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
75 802 112 826
85 810 101 826
2 B3
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
