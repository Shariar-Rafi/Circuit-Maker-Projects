CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
740 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
28
13 Logic Switch~
5 1225 276 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44852.3 0
0
13 Logic Switch~
5 1284 555 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44852.3 0
0
13 Logic Switch~
5 307 907 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90051e-315 0
0
13 Logic Switch~
5 279 421 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90051e-315 0
0
12 Hex Display~
7 1656 51 0 18 19
10 7 6 5 23 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
8157 0 0
2
44852.3 0
0
5 4030~
219 1841 240 0 3 22
0 4 3 5
0
0 0 624 90
4 4030
-7 -24 21 -16
3 U6C
26 -3 47 5
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 6 0
1 U
5572 0 0
2
44852.3 0
0
5 4030~
219 1660 236 0 3 22
0 4 2 6
0
0 0 624 90
4 4030
-7 -24 21 -16
3 U6B
26 -3 47 5
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
8901 0 0
2
44852.3 0
0
5 4030~
219 1469 233 0 3 22
0 4 10 7
0
0 0 624 90
4 4030
-7 -24 21 -16
3 U6A
26 -3 47 5
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
7361 0 0
2
44852.3 0
0
6 74112~
219 1438 451 0 7 32
0 8 8 9 8 8 24 10
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U5A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 5 0
1 U
4747 0 0
2
44852.3 4
0
6 74112~
219 1592 454 0 7 32
0 8 8 10 8 8 25 2
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U4B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 4 0
1 U
972 0 0
2
44852.3 3
0
6 74112~
219 1772 455 0 7 32
0 8 8 2 8 8 26 3
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U4A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
3472 0 0
2
44852.3 2
0
7 Pulser~
4 1193 432 0 10 12
0 27 9 28 9 0 0 5 5 1
8
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9998 0 0
2
44852.3 1
0
6 74112~
219 461 803 0 7 32
0 16 16 17 16 16 14 15
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 3 0
1 U
3536 0 0
2
5.90051e-315 5.38788e-315
0
6 74112~
219 615 806 0 7 32
0 16 16 14 16 16 13 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 3 0
1 U
4597 0 0
2
5.90051e-315 5.37752e-315
0
6 74112~
219 795 807 0 7 32
0 16 16 13 16 16 29 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3835 0 0
2
5.90051e-315 5.36716e-315
0
7 Pulser~
4 216 784 0 10 12
0 30 17 31 17 0 0 5 5 1
8
0
0 0 4656 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3670 0 0
2
5.90051e-315 5.3568e-315
0
14 Logic Display~
6 525 624 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.90051e-315 5.34643e-315
0
14 Logic Display~
6 706 624 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.90051e-315 5.32571e-315
0
14 Logic Display~
6 926 626 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.90051e-315 5.30499e-315
0
12 Hex Display~
7 344 597 0 18 19
10 15 12 11 32 0 0 0 0 0
0 1 1 1 0 0 0 0 7
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3108 0 0
2
5.90051e-315 5.26354e-315
0
12 Hex Display~
7 316 111 0 18 19
10 20 19 18 33 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
4299 0 0
2
5.90051e-315 0
0
14 Logic Display~
6 898 140 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.90051e-315 0
0
14 Logic Display~
6 678 138 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.90051e-315 0
0
14 Logic Display~
6 497 138 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
5.90051e-315 0
0
7 Pulser~
4 188 298 0 10 12
0 34 22 35 22 0 0 5 5 1
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9172 0 0
2
5.90051e-315 0
0
6 74112~
219 767 321 0 7 32
0 21 21 19 21 21 36 18
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
7100 0 0
2
5.90051e-315 0
0
6 74112~
219 587 320 0 7 32
0 21 21 20 21 21 37 19
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
3820 0 0
2
5.90051e-315 0
0
6 74112~
219 433 317 0 7 32
0 21 21 22 21 21 38 20
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
7678 0 0
2
5.90051e-315 0
0
72
0 0 2 0 0 8192 0 0 0 16 3 4
1684 323
1677 323
1677 284
1672 284
2 0 3 0 0 8192 0 6 0 0 15 3
1853 259
1853 305
1903 305
2 0 2 0 0 0 0 7 0 0 16 3
1672 255
1672 294
1683 294
1 0 4 0 0 4096 0 7 0 0 6 2
1654 255
1654 276
1 0 4 0 0 4096 0 8 0 0 6 2
1463 252
1463 276
1 1 4 0 0 4224 0 1 6 0 0 3
1237 276
1835 276
1835 259
3 3 5 0 0 8320 0 6 5 0 0 4
1844 210
1844 93
1653 93
1653 75
3 2 6 0 0 4224 0 7 5 0 0 4
1663 206
1663 88
1659 88
1659 75
3 1 7 0 0 8320 0 8 5 0 0 4
1472 203
1472 83
1665 83
1665 75
1 0 8 0 0 12288 0 11 0 0 25 4
1772 392
1772 383
1737 383
1737 555
1 0 8 0 0 0 0 10 0 0 25 4
1592 391
1592 387
1665 387
1665 555
1 0 8 0 0 0 0 9 0 0 25 4
1438 388
1438 384
1488 384
1488 555
0 3 9 0 0 4224 0 0 9 14 0 2
1227 424
1408 424
4 2 9 0 0 0 0 12 12 0 0 6
1223 432
1227 432
1227 409
1155 409
1155 432
1163 432
7 1 3 0 0 8320 0 11 0 0 0 3
1796 419
1903 419
1903 292
0 1 2 0 0 4224 0 0 0 18 0 4
1684 418
1684 298
1683 298
1683 290
0 2 10 0 0 4224 0 0 8 19 0 4
1502 415
1502 290
1481 290
1481 252
7 3 2 0 0 0 0 10 11 0 0 4
1616 418
1729 418
1729 428
1742 428
7 3 10 0 0 0 0 9 10 0 0 4
1462 415
1549 415
1549 427
1562 427
0 0 8 0 0 0 0 0 0 26 25 4
1740 437
1740 388
1733 388
1733 555
0 0 8 0 0 0 0 0 0 27 25 4
1563 436
1563 387
1557 387
1557 555
0 0 8 0 0 0 0 0 0 28 25 4
1409 433
1409 384
1403 384
1403 555
0 5 8 0 0 0 0 0 9 25 0 2
1438 555
1438 463
5 0 8 0 0 0 0 10 0 0 25 2
1592 466
1592 555
1 5 8 0 0 4224 0 2 11 0 0 3
1296 555
1772 555
1772 467
2 4 8 0 0 0 0 11 11 0 0 4
1748 419
1734 419
1734 437
1748 437
2 4 8 0 0 0 0 10 10 0 0 4
1568 418
1554 418
1554 436
1568 436
2 4 8 0 0 0 0 9 9 0 0 4
1414 415
1400 415
1400 433
1414 433
3 0 11 0 0 8320 0 20 0 0 30 3
341 621
341 719
926 719
7 1 11 0 0 0 0 15 19 0 0 3
819 771
926 771
926 644
7 0 12 0 0 8192 0 14 0 0 40 4
639 770
702 770
702 677
707 677
6 3 13 0 0 4224 0 14 15 0 0 4
645 788
752 788
752 780
765 780
6 3 14 0 0 4224 0 13 14 0 0 4
491 785
572 785
572 779
585 779
1 0 15 0 0 8320 0 20 0 0 41 3
353 621
353 660
525 660
1 0 16 0 0 12288 0 15 0 0 47 4
795 744
795 735
760 735
760 907
1 0 16 0 0 0 0 14 0 0 47 4
615 743
615 739
688 739
688 907
1 0 16 0 0 0 0 13 0 0 47 4
461 740
461 736
511 736
511 907
0 3 17 0 0 4224 0 0 13 39 0 2
250 776
431 776
4 2 17 0 0 0 0 16 16 0 0 6
246 784
250 784
250 761
178 761
178 784
186 784
1 2 12 0 0 16512 0 18 20 0 0 6
706 642
706 650
707 650
707 677
347 677
347 621
1 7 15 0 0 0 0 17 13 0 0 3
525 642
525 767
485 767
0 0 16 0 0 0 0 0 0 48 47 4
763 789
763 740
756 740
756 907
0 0 16 0 0 0 0 0 0 49 47 4
586 788
586 739
580 739
580 907
0 0 16 0 0 0 0 0 0 50 47 4
432 785
432 736
426 736
426 907
0 5 16 0 0 0 0 0 13 47 0 2
461 907
461 815
5 0 16 0 0 0 0 14 0 0 47 2
615 818
615 907
1 5 16 0 0 4224 0 3 15 0 0 3
319 907
795 907
795 819
2 4 16 0 0 0 0 15 15 0 0 4
771 771
757 771
757 789
771 789
2 4 16 0 0 0 0 14 14 0 0 4
591 770
577 770
577 788
591 788
2 4 16 0 0 0 0 13 13 0 0 4
437 767
423 767
423 785
437 785
3 0 18 0 0 8320 0 21 0 0 59 3
313 135
313 232
898 232
2 0 19 0 0 8320 0 21 0 0 60 3
319 135
319 191
679 191
1 0 20 0 0 8320 0 21 0 0 61 3
325 135
325 174
497 174
1 0 21 0 0 12288 0 26 0 0 69 4
767 258
767 249
732 249
732 421
1 0 21 0 0 0 0 27 0 0 69 4
587 257
587 253
660 253
660 421
1 0 21 0 0 0 0 28 0 0 69 4
433 254
433 250
483 250
483 421
0 3 22 0 0 4224 0 0 28 58 0 2
222 290
403 290
4 2 22 0 0 0 0 25 25 0 0 6
218 298
222 298
222 275
150 275
150 298
158 298
7 1 18 0 0 0 0 26 22 0 0 3
791 285
898 285
898 158
0 1 19 0 0 0 0 0 23 62 0 4
679 284
679 164
678 164
678 156
0 1 20 0 0 0 0 0 24 63 0 2
497 281
497 156
7 3 19 0 0 0 0 27 26 0 0 4
611 284
724 284
724 294
737 294
7 3 20 0 0 0 0 28 27 0 0 4
457 281
544 281
544 293
557 293
0 0 21 0 0 0 0 0 0 70 69 4
735 303
735 254
728 254
728 421
0 0 21 0 0 0 0 0 0 71 69 4
558 302
558 253
552 253
552 421
0 0 21 0 0 0 0 0 0 72 69 4
404 299
404 250
398 250
398 421
0 5 21 0 0 0 0 0 28 69 0 2
433 421
433 329
5 0 21 0 0 0 0 27 0 0 69 2
587 332
587 421
1 5 21 0 0 4224 0 4 26 0 0 3
291 421
767 421
767 333
2 4 21 0 0 0 0 26 26 0 0 4
743 285
729 285
729 303
743 303
2 4 21 0 0 0 0 27 27 0 0 4
563 284
549 284
549 302
563 302
2 4 21 0 0 0 0 28 28 0 0 4
409 281
395 281
395 299
409 299
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
1888 24 2013 48
1898 32 2002 48
13 mod 8 up-down
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
645 31 794 55
655 39 783 55
16 MOD 8 Up Counter
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
673 518 838 542
683 526 827 542
18 MOD 8 down counter
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
