CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
216 93 1364 691
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
426 213 567 334
9437202 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 143 266 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90047e-315 5.38788e-315
0
13 Logic Switch~
5 146 307 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V19
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90047e-315 5.37752e-315
0
13 Logic Switch~
5 193 130 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V20
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90047e-315 5.36716e-315
0
13 Logic Switch~
5 200 530 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -15 8 -7
3 V21
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90047e-315 5.3568e-315
0
13 Logic Switch~
5 235 442 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -15 8 -7
3 V22
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90047e-315 5.34643e-315
0
13 Logic Switch~
5 547 151 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V23
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90047e-315 5.32571e-315
0
13 Logic Switch~
5 607 148 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V24
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90047e-315 5.30499e-315
0
13 Logic Switch~
5 656 150 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V25
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.90047e-315 5.26354e-315
0
13 Logic Switch~
5 704 149 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V26
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.90047e-315 0
0
7 74LS194
49 472 334 0 14 29
0 15 13 14 12 11 10 2 3 4
5 6 7 8 9
0
0 0 4848 0
6 74F194
-21 -60 21 -52
3 U16
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
972 0 0
2
5.90047e-315 5.41896e-315
0
7 Pulser~
4 286 375 0 10 12
0 15 16 15 17 0 0 5 5 5
8
0
0 0 4656 0
0
3 V17
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3472 0 0
2
5.90047e-315 5.41378e-315
0
14 Logic Display~
6 885 264 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.90047e-315 5.4086e-315
0
14 Logic Display~
6 917 262 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
5.90047e-315 5.40342e-315
0
14 Logic Display~
6 950 265 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
5.90047e-315 5.39824e-315
0
14 Logic Display~
6 984 264 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-10 -28 11 -20
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
5.90047e-315 5.39306e-315
0
15
7 1 2 0 0 8320 0 10 6 0 0 4
504 298
568 298
568 151
559 151
8 1 3 0 0 8320 0 10 7 0 0 4
504 307
628 307
628 148
619 148
9 1 4 0 0 4224 0 10 8 0 0 4
504 316
677 316
677 150
668 150
10 1 5 0 0 4224 0 10 9 0 0 4
504 325
725 325
725 149
716 149
11 1 6 0 0 4224 0 10 12 0 0 3
504 343
885 343
885 282
12 1 7 0 0 4224 0 10 13 0 0 3
504 352
917 352
917 280
13 1 8 0 0 4224 0 10 14 0 0 3
504 361
950 361
950 283
14 1 9 0 0 4224 0 10 15 0 0 3
504 370
984 370
984 282
1 6 10 0 0 4224 0 5 10 0 0 4
247 442
426 442
426 370
434 370
1 5 11 0 0 4224 0 4 10 0 0 4
212 530
421 530
421 352
440 352
1 4 12 0 0 8320 0 3 10 0 0 4
205 130
411 130
411 343
440 343
1 2 13 0 0 4224 0 2 10 0 0 4
158 307
416 307
416 316
440 316
1 3 14 0 0 8320 0 1 10 0 0 5
155 266
155 322
421 322
421 325
440 325
1 0 15 0 0 12288 0 11 0 0 15 5
262 366
252 366
252 352
345 352
345 366
3 1 15 0 0 4224 0 11 10 0 0 4
310 366
426 366
426 298
440 298
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
410 8 599 32
420 16 588 32
21 4 bit universal shift
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
174 75 219 99
184 83 208 99
3 DSR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
179 538 224 562
189 546 213 562
3 DSL
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
843 216 888 240
853 224 877 240
3 MSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1010 222 1055 246
1020 230 1044 246
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
727 95 772 119
737 103 761 119
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
507 97 552 121
517 105 541 121
3 MSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
87 296 124 320
97 304 113 320
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
87 253 124 277
97 261 113 277
2 S0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
