CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 200 403 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
317 0 0
2
44851.9 0
0
13 Logic Switch~
5 198 229 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3108 0 0
2
44851.9 0
0
14 Logic Display~
6 1122 107 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4299 0 0
2
44851.9 0
0
14 Logic Display~
6 1029 109 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9672 0 0
2
44851.9 0
0
7 Pulser~
4 113 305 0 10 12
0 9 6 10 6 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7876 0 0
2
44851.9 0
0
5 7412~
219 333 394 0 4 22
0 6 5 3 7
0
0 0 624 0
6 74LS12
-14 -24 28 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 2 2 0
1 U
6369 0 0
2
44851.9 0
0
5 7412~
219 333 232 0 4 22
0 2 4 6 8
0
0 0 624 0
6 74LS12
-14 -24 28 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 1 2 0
1 U
9172 0 0
2
44851.9 0
0
5 4011~
219 758 391 0 3 22
0 3 7 2
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 1 0
1 U
7100 0 0
2
44851.9 0
0
5 4011~
219 757 230 0 3 22
0 8 2 3
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 1 0
1 U
3820 0 0
2
44851.9 0
0
14
0 0 2 0 0 8192 0 0 0 11 3 4
723 239
723 371
865 371
865 391
1 0 2 0 0 12416 0 7 0 0 3 5
309 223
295 223
295 414
800 414
800 391
3 1 2 0 0 0 0 8 3 0 0 3
785 391
1122 391
1122 125
0 1 3 0 0 4096 0 0 4 5 0 3
792 230
1029 230
1029 127
3 3 3 0 0 12416 0 6 9 0 0 6
309 403
305 403
305 210
792 210
792 230
784 230
1 2 4 0 0 4224 0 2 7 0 0 4
210 229
301 229
301 232
309 232
1 2 5 0 0 4224 0 1 6 0 0 4
212 403
301 403
301 394
309 394
0 0 6 0 0 4224 0 0 0 9 10 2
151 293
301 293
2 4 6 0 0 0 0 5 5 0 0 6
83 305
79 305
79 282
151 282
151 305
143 305
1 3 6 0 0 0 0 6 7 0 0 4
309 385
301 385
301 241
309 241
2 0 2 0 0 128 0 9 0 0 0 2
733 239
720 239
0 1 3 0 0 128 0 0 8 4 0 5
856 230
856 250
729 250
729 382
734 382
4 2 7 0 0 4224 0 6 8 0 0 4
360 394
726 394
726 400
734 400
4 1 8 0 0 4224 0 7 9 0 0 4
360 232
725 232
725 221
733 221
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 26
384 36 501 80
394 44 490 76
26 JK Flip Flop
____________
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
