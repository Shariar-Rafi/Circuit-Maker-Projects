CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 820 30 100 10
216 93 1364 691
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.390953 0.500000
426 213 567 334
9437202 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 154 629 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90046e-315 5.39306e-315
0
13 Logic Switch~
5 130 841 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90046e-315 5.38788e-315
0
13 Logic Switch~
5 115 587 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.90046e-315 5.37752e-315
0
13 Logic Switch~
5 101 125 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90046e-315 5.30499e-315
0
13 Logic Switch~
5 112 378 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90046e-315 5.26354e-315
0
13 Logic Switch~
5 140 167 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90046e-315 0
0
12 Hex Display~
7 698 502 0 18 19
10 11 10 9 40 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
8901 0 0
2
5.90046e-315 0
0
12 Hex Display~
7 697 37 0 18 19
10 15 14 13 41 0 0 0 0 0
0 1 1 1 0 0 0 0 7
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
7361 0 0
2
5.90046e-315 0
0
14 Logic Display~
6 622 512 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.90046e-315 5.36716e-315
0
14 Logic Display~
6 468 515 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.90046e-315 5.3568e-315
0
14 Logic Display~
6 321 511 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.90046e-315 5.34643e-315
0
6 74112~
219 529 722 0 7 32
0 18 12 16 12 19 42 9
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 3 0
1 U
9998 0 0
2
5.90046e-315 5.32571e-315
0
6 74112~
219 405 722 0 7 32
0 18 12 17 12 19 16 10
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 3 0
1 U
3536 0 0
2
5.90046e-315 5.30499e-315
0
6 74112~
219 264 715 0 7 32
0 18 12 20 12 19 17 11
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 2 0
1 U
4597 0 0
2
5.90046e-315 5.26354e-315
0
7 Pulser~
4 123 697 0 10 12
0 20 43 20 44 0 0 10 10 1
8
0
0 0 4640 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3835 0 0
2
5.90046e-315 0
0
7 Pulser~
4 109 235 0 10 12
0 24 45 24 46 0 0 10 10 1
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3670 0 0
2
5.90046e-315 5.39306e-315
0
6 74112~
219 250 253 0 7 32
0 22 21 24 21 23 47 15
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
5616 0 0
2
5.90046e-315 5.38788e-315
0
6 74112~
219 391 260 0 7 32
0 22 21 15 21 23 48 14
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
9323 0 0
2
5.90046e-315 5.37752e-315
0
6 74112~
219 515 260 0 7 32
0 22 21 14 21 23 49 13
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
317 0 0
2
5.90046e-315 5.36716e-315
0
14 Logic Display~
6 307 49 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.90046e-315 5.3568e-315
0
14 Logic Display~
6 454 53 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
5.90046e-315 5.34643e-315
0
14 Logic Display~
6 608 50 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.90046e-315 5.32571e-315
0
44
0 3 9 0 0 4096 0 0 7 4 0 3
622 561
695 561
695 526
2 0 10 0 0 8320 0 7 0 0 5 3
701 526
701 568
468 568
1 0 11 0 0 8320 0 7 0 0 6 3
707 526
707 575
321 575
7 1 9 0 0 8320 0 12 9 0 0 3
553 686
622 686
622 530
7 1 10 0 0 0 0 13 10 0 0 3
429 686
468 686
468 533
7 1 11 0 0 0 0 14 11 0 0 3
288 679
321 679
321 529
4 0 12 0 0 8192 0 12 0 0 17 3
505 704
482 704
482 629
4 0 12 0 0 0 0 13 0 0 17 3
381 704
346 704
346 629
2 0 12 0 0 0 0 13 0 0 17 3
381 686
329 686
329 629
4 0 12 0 0 0 0 14 0 0 17 3
240 697
186 697
186 629
2 0 12 0 0 0 0 14 0 0 17 3
240 679
178 679
178 629
1 3 13 0 0 8192 0 22 8 0 0 4
608 68
608 72
694 72
694 61
2 0 14 0 0 8320 0 8 0 0 35 3
700 61
700 77
454 77
1 0 15 0 0 8320 0 8 0 0 36 3
706 61
706 93
307 93
6 3 16 0 0 4224 0 13 12 0 0 4
435 704
491 704
491 695
499 695
6 3 17 0 0 4224 0 14 13 0 0 4
294 697
362 697
362 695
375 695
1 2 12 0 0 4224 0 1 12 0 0 4
166 629
491 629
491 686
505 686
1 0 18 0 0 4096 0 13 0 0 23 2
405 659
405 587
1 0 18 0 0 0 0 14 0 0 23 2
264 652
264 587
5 0 19 0 0 4096 0 14 0 0 22 2
264 727
264 840
5 0 19 0 0 0 0 13 0 0 22 2
405 734
405 840
1 5 19 0 0 12416 0 2 12 0 0 5
142 841
264 841
264 840
529 840
529 734
1 1 18 0 0 4224 0 3 12 0 0 3
127 587
529 587
529 659
0 3 20 0 0 4224 0 0 14 25 0 2
161 688
234 688
1 3 20 0 0 0 0 15 15 0 0 6
99 688
89 688
89 674
161 674
161 688
147 688
4 0 21 0 0 8192 0 19 0 0 31 3
491 242
481 242
481 224
4 0 21 0 0 0 0 17 0 0 30 3
226 235
216 235
216 217
4 0 21 0 0 0 0 18 0 0 29 3
367 242
355 242
355 224
2 0 21 0 0 8192 0 18 0 0 31 3
367 224
346 224
346 167
2 0 21 0 0 0 0 17 0 0 31 3
226 217
216 217
216 167
1 2 21 0 0 4224 0 6 19 0 0 4
152 167
477 167
477 224
491 224
0 3 14 0 0 0 0 0 19 35 0 3
431 224
431 233
485 233
3 0 15 0 0 0 0 18 0 0 36 3
361 233
287 233
287 217
7 1 13 0 0 8320 0 19 22 0 0 3
539 224
608 224
608 68
7 1 14 0 0 0 0 18 21 0 0 3
415 224
454 224
454 71
7 1 15 0 0 0 0 17 20 0 0 3
274 217
307 217
307 67
1 0 22 0 0 4096 0 18 0 0 42 2
391 197
391 125
1 0 22 0 0 0 0 17 0 0 42 2
250 190
250 125
5 0 23 0 0 4096 0 17 0 0 41 2
250 265
250 378
5 0 23 0 0 0 0 18 0 0 41 2
391 272
391 378
1 5 23 0 0 4224 0 5 19 0 0 3
124 378
515 378
515 272
1 1 22 0 0 4224 0 4 19 0 0 3
113 125
515 125
515 197
0 3 24 0 0 4224 0 0 17 44 0 2
147 226
220 226
1 3 24 0 0 0 0 16 16 0 0 6
85 226
75 226
75 212
147 212
147 226
133 226
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 52
6 3 219 47
12 7 212 39
52 JK up counter with mod 8:
-------------------------
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 56
7 455 236 499
13 459 229 491
56 JK down counter with mod 8:
---------------------------
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
898 1 967 85
904 5 960 69
27 Lab 
Group
NO-5
_______
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
