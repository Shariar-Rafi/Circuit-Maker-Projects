CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 538 475 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44829.5 0
0
13 Logic Switch~
5 413 481 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44829.5 1
0
13 Logic Switch~
5 248 483 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44829.5 2
0
13 Logic Switch~
5 98 426 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
44829.5 3
0
13 Logic Switch~
5 85 142 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
44829.5 4
0
13 Logic Switch~
5 127 486 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-8 -17 6 -9
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
44829.5 5
0
5 4013~
219 575 282 0 6 22
0 12 9 6 5 13 7
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U8B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 4 0
1 U
8901 0 0
2
44829.5 6
0
5 4013~
219 476 282 0 6 22
0 12 10 6 5 14 8
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U8A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 4 0
1 U
7361 0 0
2
44829.5 7
0
5 4013~
219 352 297 0 6 22
0 12 4 6 5 15 2
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U7B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 3 0
1 U
4747 0 0
2
44829.5 8
0
5 4013~
219 210 288 0 6 22
0 12 11 6 5 16 3
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U7A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 3 0
1 U
972 0 0
2
44829.5 9
0
14 Logic Display~
6 884 118 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
44829.5 10
0
14 Logic Display~
6 847 120 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
44829.5 11
0
14 Logic Display~
6 808 122 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
44829.5 12
0
14 Logic Display~
6 763 111 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
44829.5 13
0
7 Pulser~
4 94 305 0 10 12
0 6 17 6 18 0 0 5 5 1
8
0
0 0 4656 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3835 0 0
2
44829.5 14
0
24
6 1 2 0 0 16512 0 9 13 0 0 6
376 261
376 219
448 219
448 174
808 174
808 140
6 1 3 0 0 12416 0 10 14 0 0 5
234 252
324 252
324 193
763 193
763 129
1 2 4 0 0 8320 0 3 9 0 0 4
260 483
315 483
315 261
328 261
4 0 5 0 0 4096 0 7 0 0 15 3
575 288
575 306
576 306
4 0 5 0 0 0 0 8 0 0 12 2
476 288
476 305
3 0 6 0 0 4096 0 9 0 0 21 3
328 279
328 274
326 274
6 1 7 0 0 4224 0 7 11 0 0 3
599 246
884 246
884 136
6 1 8 0 0 12416 0 8 12 0 0 7
500 246
543 246
543 213
834 213
834 146
847 146
847 138
1 2 9 0 0 8320 0 1 7 0 0 6
550 475
555 475
555 306
547 306
547 246
551 246
1 2 10 0 0 8320 0 2 8 0 0 4
425 481
444 481
444 246
452 246
1 2 11 0 0 8320 0 6 10 0 0 4
139 486
178 486
178 252
186 252
0 0 5 0 0 4096 0 0 0 0 15 4
476 302
476 421
477 421
477 426
4 0 5 0 0 0 0 9 0 0 15 4
352 303
352 411
355 411
355 426
0 4 5 0 0 4096 0 0 10 15 0 2
210 426
210 294
1 0 5 0 0 4224 0 4 0 0 0 3
110 426
576 426
576 302
1 0 12 0 0 4096 0 8 0 0 19 2
476 225
476 142
1 0 12 0 0 0 0 9 0 0 19 4
352 240
352 157
355 157
355 142
1 0 12 0 0 4096 0 10 0 0 19 2
210 231
210 142
1 1 12 0 0 4224 0 5 7 0 0 4
97 142
576 142
576 225
575 225
0 3 6 0 0 4096 0 0 8 24 0 3
432 313
432 264
452 264
0 0 6 0 0 0 0 0 0 24 0 3
320 313
320 274
331 274
0 3 6 0 0 0 0 0 10 24 0 3
174 296
174 270
186 270
1 0 6 0 0 12288 0 15 0 0 24 5
70 296
60 296
60 282
149 282
149 296
3 3 6 0 0 12416 0 15 7 0 0 6
118 296
182 296
182 313
544 313
544 264
551 264
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
929 2 1078 26
939 10 1067 26
16 (Input = Output)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
359 162 412 186
369 170 401 186
4 PIPO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
311 56 364 80
321 64 353 80
4 PIPO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
117 501 146 525
123 505 139 521
2 P3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
239 502 268 526
245 506 261 522
2 P2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
399 493 428 517
405 497 421 513
2 P3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
531 494 560 538
537 498 553 530
2 P4
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
