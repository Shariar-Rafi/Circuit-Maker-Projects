CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 171 118 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44852 0
0
14 Logic Display~
6 887 280 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
391 0 0
2
44852 0
0
14 Logic Display~
6 884 164 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3124 0 0
2
44852 0
0
7 Pulser~
4 84 228 0 10 12
0 9 7 10 7 0 0 5 5 4
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3421 0 0
2
44852 0
0
9 Inverter~
13 253 313 0 2 22
0 6 8
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
8157 0 0
2
44852 0
0
10 2-In NAND~
219 619 300 0 3 22
0 2 5 3
0
0 0 624 0
5 74F37
-10 -24 25 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
5572 0 0
2
44852 0
0
10 2-In NAND~
219 619 190 0 3 22
0 4 3 2
0
0 0 624 0
5 74F37
-10 -24 25 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
8901 0 0
2
44852 0
0
10 2-In NAND~
219 364 302 0 3 22
0 7 8 5
0
0 0 624 0
5 74F37
-10 -24 25 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7361 0 0
2
44852 0
0
10 2-In NAND~
219 361 192 0 3 22
0 6 7 4
0
0 0 624 0
5 74F37
-10 -24 25 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4747 0 0
2
44852 0
0
13
1 0 2 0 0 8192 0 6 0 0 8 5
595 291
581 291
581 170
687 170
687 190
2 0 3 0 0 8192 0 7 0 0 9 5
595 199
591 199
591 320
691 320
691 300
3 1 4 0 0 4224 0 9 7 0 0 4
388 192
587 192
587 181
595 181
3 2 5 0 0 4224 0 8 6 0 0 4
391 302
587 302
587 309
595 309
0 1 6 0 0 4096 0 0 9 6 0 2
230 183
337 183
0 0 6 0 0 0 0 0 0 7 0 2
230 118
230 183
1 1 6 0 0 8320 0 1 5 0 0 4
183 118
230 118
230 313
238 313
3 1 2 0 0 4224 0 7 3 0 0 3
646 190
884 190
884 182
3 1 3 0 0 4240 0 6 2 0 0 3
646 300
887 300
887 298
0 0 7 0 0 4224 0 0 0 12 11 2
122 218
329 218
1 2 7 0 0 0 0 8 9 0 0 4
340 293
329 293
329 201
337 201
2 4 7 0 0 0 0 4 4 0 0 6
54 228
50 228
50 205
122 205
122 228
114 228
2 2 8 0 0 4224 0 5 8 0 0 4
274 313
332 313
332 311
340 311
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
375 13 484 37
385 21 473 37
11 D Flip Flop
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
