CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
261 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
429 176 542 273
9437202 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 103 312 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-8 -16 6 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44789.9 3
0
13 Logic Switch~
5 104 360 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
44789.9 2
0
13 Logic Switch~
5 101 184 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
44789.9 0
0
13 Logic Switch~
5 100 132 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
44789.9 0
0
13 Logic Switch~
5 99 84 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-8 -16 6 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
44789.9 0
0
9 2-In XOR~
219 207 330 0 3 22
0 10 9 3
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
5572 0 0
2
44789.9 7
0
9 2-In XOR~
219 400 332 0 3 22
0 3 2 5
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
8901 0 0
2
44789.9 6
0
9 2-In AND~
219 208 487 0 3 22
0 10 9 7
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
7361 0 0
2
44789.9 5
0
8 2-In OR~
219 497 470 0 3 22
0 8 7 4
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
4747 0 0
2
44789.9 4
0
9 2-In AND~
219 384 445 0 3 22
0 2 3 8
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
972 0 0
2
44789.9 0
0
14 Logic Display~
6 669 221 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
44789.9 0
0
14 Logic Display~
6 652 158 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
44789.9 0
0
14 Logic Display~
6 637 97 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
44789.9 0
0
9 2-In AND~
219 361 228 0 3 22
0 14 13 12
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
4597 0 0
2
44789.9 0
0
8 2-In OR~
219 493 242 0 3 22
0 12 11 2
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3835 0 0
2
44789.9 0
0
9 2-In AND~
219 204 259 0 3 22
0 16 15 11
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3670 0 0
2
44789.9 0
0
9 2-In XOR~
219 396 104 0 3 22
0 14 13 6
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
5616 0 0
2
44789.9 0
0
9 2-In XOR~
219 203 102 0 3 22
0 16 15 14
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9323 0 0
2
44789.9 0
0
23
0 1 2 0 0 4096 0 0 10 6 0 5
397 352
397 426
352 426
352 436
360 436
0 2 3 0 0 4096 0 0 10 11 0 3
266 330
266 454
360 454
3 1 4 0 0 8320 0 9 11 0 0 3
530 470
669 470
669 239
3 1 5 0 0 4224 0 7 12 0 0 3
433 332
652 332
652 176
3 1 6 0 0 8336 0 17 13 0 0 4
429 104
429 125
637 125
637 115
3 2 2 0 0 12416 0 15 7 0 0 6
526 242
530 242
530 352
376 352
376 341
384 341
3 2 7 0 0 4224 0 8 9 0 0 4
229 487
465 487
465 479
484 479
3 1 8 0 0 4224 0 10 9 0 0 4
405 445
462 445
462 461
484 461
0 2 9 0 0 4224 0 0 8 12 0 3
139 360
139 496
184 496
0 1 10 0 0 4224 0 0 8 13 0 3
163 312
163 478
184 478
3 1 3 0 0 4224 0 6 7 0 0 4
240 330
376 330
376 323
384 323
1 2 9 0 0 0 0 2 6 0 0 4
116 360
183 360
183 339
191 339
1 1 10 0 0 0 0 1 6 0 0 4
115 312
183 312
183 321
191 321
3 2 11 0 0 4224 0 16 15 0 0 4
225 259
461 259
461 251
480 251
3 1 12 0 0 4224 0 14 15 0 0 4
382 228
458 228
458 233
480 233
0 2 13 0 0 4096 0 0 14 20 0 3
304 184
304 237
337 237
1 0 14 0 0 8192 0 14 0 0 21 3
337 219
329 219
329 102
0 2 15 0 0 4224 0 0 16 22 0 3
135 132
135 268
180 268
0 1 16 0 0 4224 0 0 16 23 0 3
159 84
159 250
180 250
1 2 13 0 0 4224 0 3 17 0 0 4
113 184
372 184
372 113
380 113
3 1 14 0 0 4224 0 18 17 0 0 4
236 102
372 102
372 95
380 95
1 2 15 0 0 0 0 4 18 0 0 4
112 132
179 132
179 111
187 111
1 1 16 0 0 0 0 5 18 0 0 4
111 84
179 84
179 93
187 93
45
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
343 329 380 353
353 337 369 353
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
359 299 396 323
369 307 385 323
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
421 303 454 327
429 311 445 327
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
523 445 548 469
531 452 539 468
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
469 476 494 500
477 484 485 500
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
466 442 491 466
474 450 482 466
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
220 462 257 486
230 470 246 486
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
164 493 201 517
174 501 190 517
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
164 454 201 478
174 462 190 478
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
339 451 376 475
349 459 365 475
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
334 418 359 442
342 426 350 442
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
405 422 434 446
415 430 423 446
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
174 345 211 369
184 353 200 369
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
232 305 257 329
240 313 248 329
1 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
170 291 195 315
178 298 186 314
1 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
465 249 490 273
473 257 481 273
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
516 218 541 242
524 226 532 242
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
464 211 489 235
472 219 480 235
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
375 207 400 231
383 215 391 231
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
325 234 350 258
333 242 341 258
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
327 196 352 220
335 204 343 220
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
165 227 190 251
173 235 181 251
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
221 235 250 259
231 243 239 259
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
163 263 192 287
173 271 181 287
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
844 86 905 110
854 94 894 110
5 Note:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
851 134 876 158
859 141 867 157
1 +
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
856 156 901 180
866 164 890 180
3 101
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
861 131 898 155
871 138 887 154
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
860 107 897 131
870 115 886 131
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
370 117 399 141
380 125 388 141
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
366 72 391 96
374 80 382 96
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
432 99 461 123
442 107 450 123
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
159 50 184 74
167 58 175 74
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
230 80 259 104
240 88 248 104
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
171 115 200 139
181 123 189 139
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
636 469 673 493
646 477 662 493
2 C2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
586 330 623 354
596 338 612 354
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
534 239 571 263
544 247 560 263
2 C1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
509 91 546 115
519 99 535 115
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
51 342 88 366
61 349 77 365
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
47 296 84 320
57 304 73 320
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
50 115 83 139
58 123 74 139
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
52 66 85 90
60 74 76 90
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
246 3 363 27
256 11 352 27
12 2 Bit Adder:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
41 169 94 193
51 177 83 193
4 C0=0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
