CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
216 93 1364 691
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
426 213 567 334
42991634 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 754 2123 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V26
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44824.4 1
0
13 Logic Switch~
5 706 2124 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V25
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44824.4 2
0
13 Logic Switch~
5 657 2122 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V24
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44824.4 3
0
13 Logic Switch~
5 597 2125 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V23
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
44824.4 4
0
13 Logic Switch~
5 285 2416 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -15 8 -7
3 V22
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
44824.4 5
0
13 Logic Switch~
5 250 2504 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -15 8 -7
3 V21
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
44824.4 6
0
13 Logic Switch~
5 243 2104 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V20
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
44824.4 7
0
13 Logic Switch~
5 196 2281 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V19
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
44824.4 8
0
13 Logic Switch~
5 193 2240 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V18
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
44824.4 9
0
13 Logic Switch~
5 117 187 0 10 11
0 58 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
44824.4 21
0
14 Logic Display~
6 1034 2238 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -28 11 -20
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
44824.4 22
0
14 Logic Display~
6 1000 2239 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
44824.4 23
0
14 Logic Display~
6 967 2236 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
44824.4 24
0
14 Logic Display~
6 935 2238 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
44824.4 25
0
7 Pulser~
4 336 2349 0 10 12
0 19 59 19 60 0 0 5 5 6
7
0
0 0 4640 0
0
3 V17
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3835 0 0
2
44824.4 26
0
7 74LS194
49 522 2308 0 14 29
0 19 17 18 16 15 14 3 4 5
6 7 8 9 10
0
0 0 4832 0
6 74F194
-21 -60 21 -52
3 U16
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
3670 0 0
2
44824.4 27
0
14 Logic Display~
6 629 64 0 1 2
10 54
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
44824.4 62
0
7 Pulser~
4 121 276 0 10 12
0 53 79 53 80 0 0 5 5 6
7
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9323 0 0
2
44824.4 63
0
12 D Flip-Flop~
219 585 239 0 4 9
0 55 53 81 54
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U4
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
317 0 0
2
44824.4 64
0
12 D Flip-Flop~
219 492 241 0 4 9
0 56 53 82 55
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U3
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3108 0 0
2
44824.4 65
0
12 D Flip-Flop~
219 390 243 0 4 9
0 57 53 83 56
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U2
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4299 0 0
2
44824.4 66
0
12 D Flip-Flop~
219 273 246 0 4 9
0 58 53 84 57
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U1
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9672 0 0
2
44824.4 67
0
25
7 1 3 0 0 8320 0 16 4 0 0 4
554 2272
618 2272
618 2125
609 2125
8 1 4 0 0 8320 0 16 3 0 0 4
554 2281
678 2281
678 2122
669 2122
9 1 5 0 0 4224 0 16 2 0 0 4
554 2290
727 2290
727 2124
718 2124
10 1 6 0 0 4224 0 16 1 0 0 4
554 2299
775 2299
775 2123
766 2123
11 1 7 0 0 4224 0 16 14 0 0 3
554 2317
935 2317
935 2256
12 1 8 0 0 4224 0 16 13 0 0 3
554 2326
967 2326
967 2254
13 1 9 0 0 4224 0 16 12 0 0 3
554 2335
1000 2335
1000 2257
14 1 10 0 0 4224 0 16 11 0 0 3
554 2344
1034 2344
1034 2256
1 6 14 0 0 4224 0 5 16 0 0 4
297 2416
476 2416
476 2344
484 2344
1 5 15 0 0 4224 0 6 16 0 0 4
262 2504
471 2504
471 2326
490 2326
1 4 16 0 0 8320 0 7 16 0 0 4
255 2104
461 2104
461 2317
490 2317
1 2 17 0 0 4224 0 8 16 0 0 4
208 2281
466 2281
466 2290
490 2290
1 3 18 0 0 8320 0 9 16 0 0 5
205 2240
205 2296
471 2296
471 2299
490 2299
1 0 19 0 0 12288 0 15 0 0 15 5
312 2340
302 2340
302 2326
395 2326
395 2340
3 1 19 0 0 4224 0 15 16 0 0 4
360 2340
476 2340
476 2272
490 2272
1 0 53 0 0 12288 0 18 0 0 21 5
97 267
87 267
87 242
166 242
166 267
4 1 54 0 0 8320 0 19 17 0 0 3
609 203
629 203
629 82
2 0 53 0 0 0 0 22 0 0 21 3
249 228
243 228
243 267
2 0 53 0 0 0 0 21 0 0 21 3
366 225
361 225
361 267
2 0 53 0 0 0 0 20 0 0 21 3
468 223
461 223
461 267
3 2 53 0 0 4224 0 18 19 0 0 4
145 267
553 267
553 221
561 221
4 1 55 0 0 4224 0 20 19 0 0 4
516 205
553 205
553 203
561 203
4 1 56 0 0 4224 0 21 20 0 0 4
414 207
460 207
460 205
468 205
4 1 57 0 0 4224 0 22 21 0 0 4
297 210
358 210
358 207
366 207
1 1 58 0 0 4224 0 10 22 0 0 4
129 187
241 187
241 210
249 210
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
460 1982 649 2006
470 1990 638 2006
21 4 bit universal shift
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
224 2049 269 2073
234 2057 258 2073
3 DSR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
229 2512 274 2536
239 2520 263 2536
3 DSL
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
893 2190 938 2214
903 2198 927 2214
3 MSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1060 2196 1105 2220
1070 2204 1094 2220
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
777 2069 822 2093
787 2077 811 2093
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
557 2071 602 2095
567 2079 591 2095
3 MSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
137 2270 174 2294
147 2278 163 2294
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
137 2227 174 2251
147 2235 163 2251
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
294 34 347 58
304 42 336 58
4 SISO
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
