CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
90 220 30 80 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
77 E:\Software (Installed and Running)\Electronics\CircuitMaker 2000 SP1\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
81
13 Logic Switch~
5 118 1002 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V12
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3608 0 0
2
5.90052e-315 0
0
13 Logic Switch~
5 151 1003 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V11
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6397 0 0
2
5.90052e-315 5.26354e-315
0
13 Logic Switch~
5 187 1004 0 10 11
0 44 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
3 V10
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3967 0 0
2
5.90052e-315 5.30499e-315
0
13 Logic Switch~
5 219 1004 0 10 11
0 62 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8621 0 0
2
5.90052e-315 5.32571e-315
0
13 Logic Switch~
5 217 901 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90052e-315 5.34643e-315
0
13 Logic Switch~
5 185 901 0 10 11
0 45 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7385 0 0
2
5.90052e-315 5.3568e-315
0
13 Logic Switch~
5 149 900 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6519 0 0
2
5.90052e-315 5.36716e-315
0
13 Logic Switch~
5 116 899 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
552 0 0
2
5.90052e-315 5.37752e-315
0
13 Logic Switch~
5 219 801 0 1 11
0 63
0
0 0 21360 90
2 0V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5551 0 0
2
5.90052e-315 5.38788e-315
0
13 Logic Switch~
5 187 801 0 1 11
0 7
0
0 0 21360 90
2 0V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8715 0 0
2
5.90052e-315 5.39306e-315
0
13 Logic Switch~
5 151 800 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9763 0 0
2
5.90052e-315 5.39824e-315
0
13 Logic Switch~
5 118 799 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8443 0 0
2
5.90052e-315 5.40342e-315
0
14 Logic Display~
6 1603 251 0 1 2
10 61
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3719 0 0
2
44859.8 0
0
14 Logic Display~
6 1579 251 0 1 2
10 43
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8671 0 0
2
44859.8 1
0
14 Logic Display~
6 1553 252 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
44859.8 2
0
14 Logic Display~
6 1524 251 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
49 0 0
2
44859.8 3
0
14 Logic Display~
6 1476 247 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6536 0 0
2
44859.8 4
0
9 2-In AND~
219 1031 479 0 3 22
0 34 33 41
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 18 0
1 U
3931 0 0
2
44859.8 5
0
9 2-In AND~
219 1031 525 0 3 22
0 42 39 40
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 18 0
1 U
4390 0 0
2
44859.8 6
0
8 2-In OR~
219 1082 488 0 3 22
0 41 40 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U11D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
3242 0 0
2
44859.8 7
0
9 2-In AND~
219 922 454 0 3 22
0 28 29 39
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
6760 0 0
2
44859.8 8
0
9 2-In XOR~
219 980 423 0 3 22
0 34 33 42
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U13D
-10 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
5760 0 0
2
44859.8 9
0
9 2-In XOR~
219 1064 432 0 3 22
0 42 39 25
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U13C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
3781 0 0
2
44859.8 10
0
8 2-In OR~
219 974 635 0 3 22
0 36 35 33
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U11C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
8545 0 0
2
44859.8 11
0
9 2-In AND~
219 923 672 0 3 22
0 8 32 35
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
9739 0 0
2
44859.8 12
0
9 2-In AND~
219 923 626 0 3 22
0 7 26 36
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
388 0 0
2
44859.8 13
0
5 4082~
219 923 574 0 5 22
0 31 8 9 32 37
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U17B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 17 0
1 U
4595 0 0
2
44859.8 14
0
5 4082~
219 923 527 0 5 22
0 31 30 9 26 38
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U17A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 17 0
1 U
3173 0 0
2
44859.8 15
0
8 3-In OR~
219 973 574 0 4 22
0 38 37 27 34
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U16A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 16 0
1 U
9261 0 0
2
44859.8 16
0
9 Inverter~
13 954 700 0 2 22
0 26 32
0
0 0 624 180
6 74LS04
-21 -19 21 -11
4 U15D
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 15 0
1 U
3494 0 0
2
44859.8 17
0
9 Inverter~
13 895 364 0 2 22
0 7 31
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U15C
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 15 0
1 U
9101 0 0
2
44859.8 18
0
9 Inverter~
13 943 365 0 2 22
0 8 30
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U15B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 15 0
1 U
358 0 0
2
44859.8 19
0
9 Inverter~
13 989 366 0 2 22
0 9 29
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U15A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 15 0
1 U
3726 0 0
2
44859.8 20
0
9 Inverter~
13 1287 366 0 2 22
0 9 11
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U8F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
999 0 0
2
44859.8 21
0
9 Inverter~
13 1241 365 0 2 22
0 8 12
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U8E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
8787 0 0
2
44859.8 22
0
9 Inverter~
13 1193 364 0 2 22
0 7 13
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U8D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 8 0
1 U
3348 0 0
2
44859.8 23
0
9 Inverter~
13 1252 700 0 2 22
0 5 14
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U8C
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 8 0
1 U
3395 0 0
2
44859.8 24
0
8 3-In OR~
219 1271 574 0 4 22
0 20 19 6 16
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U1C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 1 0
1 U
7740 0 0
2
44859.8 25
0
5 4082~
219 1221 527 0 5 22
0 13 12 9 5 20
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U14B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 14 0
1 U
6480 0 0
2
44859.8 26
0
5 4082~
219 1221 574 0 5 22
0 13 8 9 14 19
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U14A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 14 0
1 U
342 0 0
2
44859.8 27
0
9 2-In AND~
219 1221 626 0 3 22
0 7 5 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
9953 0 0
2
44859.8 28
0
9 2-In AND~
219 1221 672 0 3 22
0 8 14 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
361 0 0
2
44859.8 29
0
8 2-In OR~
219 1272 635 0 3 22
0 18 17 15
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U11B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
3343 0 0
2
44859.8 30
0
9 2-In XOR~
219 1362 432 0 3 22
0 24 21 3
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U13B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
7923 0 0
2
44859.8 31
0
9 2-In XOR~
219 1278 423 0 3 22
0 16 15 24
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U13A
-10 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
6174 0 0
2
44859.8 32
0
9 2-In AND~
219 1220 454 0 3 22
0 10 11 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
6692 0 0
2
44859.8 33
0
8 2-In OR~
219 1380 488 0 3 22
0 23 22 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U11A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
8790 0 0
2
44859.8 34
0
9 2-In AND~
219 1329 525 0 3 22
0 24 21 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
4595 0 0
2
44859.8 35
0
9 2-In AND~
219 1329 479 0 3 22
0 16 15 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
667 0 0
2
44859.8 36
0
9 2-In AND~
219 733 479 0 3 22
0 52 51 59
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
8743 0 0
2
44859.8 37
0
9 2-In AND~
219 733 525 0 3 22
0 60 57 58
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
8298 0 0
2
44859.8 38
0
8 2-In OR~
219 784 488 0 3 22
0 59 58 28
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
313 0 0
2
44859.8 39
0
9 2-In AND~
219 624 454 0 3 22
0 46 47 57
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
7548 0 0
2
44859.8 40
0
9 2-In XOR~
219 682 423 0 3 22
0 52 51 60
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6D
-7 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
8973 0 0
2
44859.8 41
0
9 2-In XOR~
219 766 432 0 3 22
0 60 57 43
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
9712 0 0
2
44859.8 42
0
8 2-In OR~
219 676 635 0 3 22
0 54 53 51
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
4518 0 0
2
44859.8 43
0
9 2-In AND~
219 625 672 0 3 22
0 8 50 53
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
5596 0 0
2
44859.8 44
0
9 2-In AND~
219 625 626 0 3 22
0 7 44 54
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
692 0 0
2
44859.8 45
0
5 4082~
219 625 574 0 5 22
0 49 8 9 50 55
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U9B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 9 0
1 U
6258 0 0
2
44859.8 46
0
5 4082~
219 625 527 0 5 22
0 49 48 9 44 56
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U9A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 9 0
1 U
5578 0 0
2
44859.8 47
0
8 3-In OR~
219 675 574 0 4 22
0 56 55 45 52
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U1B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 1 0
1 U
8709 0 0
2
44859.8 48
0
9 Inverter~
13 656 700 0 2 22
0 44 50
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U8B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
9131 0 0
2
44859.8 49
0
9 Inverter~
13 597 364 0 2 22
0 7 49
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U8A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
3645 0 0
2
44859.8 50
0
9 Inverter~
13 645 365 0 2 22
0 8 48
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U7F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 7 0
1 U
7613 0 0
2
44859.8 51
0
9 Inverter~
13 691 366 0 2 22
0 9 47
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U7E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 7 0
1 U
9467 0 0
2
44859.8 52
0
9 Inverter~
13 393 366 0 2 22
0 9 64
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U7D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 7 0
1 U
3932 0 0
2
5.90052e-315 5.4086e-315
0
9 Inverter~
13 347 365 0 2 22
0 8 65
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U7C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 7 0
1 U
5288 0 0
2
5.90052e-315 5.41378e-315
0
9 Inverter~
13 299 364 0 2 22
0 7 66
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U7B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 7 0
1 U
4934 0 0
2
5.90052e-315 5.41896e-315
0
9 Inverter~
13 358 700 0 2 22
0 62 67
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U7A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
5987 0 0
2
5.90052e-315 5.42414e-315
0
8 3-In OR~
219 377 574 0 4 22
0 73 72 2 69
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 1 0
1 U
7737 0 0
2
44859.8 53
0
5 4082~
219 327 527 0 5 22
0 66 65 9 62 73
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
4200 0 0
2
44859.8 54
0
5 4082~
219 327 574 0 5 22
0 66 8 9 67 72
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
5780 0 0
2
44859.8 55
0
9 2-In AND~
219 327 626 0 3 22
0 7 62 71
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6490 0 0
2
44859.8 56
0
9 2-In AND~
219 327 672 0 3 22
0 8 67 70
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8663 0 0
2
44859.8 57
0
8 2-In OR~
219 378 635 0 3 22
0 71 70 68
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
318 0 0
2
44859.8 58
0
9 2-In XOR~
219 468 432 0 3 22
0 77 74 61
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
348 0 0
2
5.90052e-315 5.42933e-315
0
9 2-In XOR~
219 384 423 0 3 22
0 69 68 77
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6A
-7 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
8551 0 0
2
5.90052e-315 5.43192e-315
0
9 2-In AND~
219 326 454 0 3 22
0 63 64 74
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7295 0 0
2
5.90052e-315 5.43451e-315
0
8 2-In OR~
219 486 488 0 3 22
0 76 75 46
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9900 0 0
2
5.90052e-315 5.4371e-315
0
9 2-In AND~
219 435 525 0 3 22
0 77 74 75
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
8725 0 0
2
5.90052e-315 5.43969e-315
0
9 2-In AND~
219 435 479 0 3 22
0 69 68 76
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
366 0 0
2
5.90052e-315 5.44228e-315
0
137
1 3 2 0 0 8320 0 5 70 0 0 9
218 888
218 866
438 866
438 737
443 737
443 599
354 599
354 583
364 583
1 3 3 0 0 4224 0 16 44 0 0 5
1524 269
1524 716
1422 716
1422 432
1395 432
1 3 4 0 0 12416 0 17 47 0 0 5
1476 265
1476 272
1441 272
1441 488
1413 488
1 0 5 0 0 8320 0 1 0 0 20 7
119 989
119 949
1319 949
1319 737
1324 737
1324 706
1306 706
1 3 6 0 0 8320 0 8 38 0 0 9
117 886
117 843
1332 843
1332 737
1337 737
1337 599
1248 599
1248 583
1258 583
1 0 7 0 0 8320 0 10 0 0 16 4
188 788
188 273
1189 273
1189 342
1 0 8 0 0 8320 0 11 0 0 14 4
152 787
152 246
1198 246
1198 337
1 0 9 0 0 12416 0 12 0 0 12 5
119 786
121 786
121 228
1207 228
1207 332
3 1 10 0 0 8320 0 20 46 0 0 9
1115 488
1143 488
1143 288
1328 288
1328 393
1264 393
1264 407
1196 407
1196 445
2 2 11 0 0 12416 0 34 46 0 0 6
1290 384
1260 384
1260 404
1192 404
1192 463
1196 463
3 0 9 0 0 0 0 39 0 0 12 2
1197 532
1171 532
1 3 9 0 0 0 0 34 40 0 0 5
1290 348
1290 332
1171 332
1171 579
1197 579
2 0 8 0 0 0 0 40 0 0 14 2
1197 570
1176 570
1 1 8 0 0 0 0 35 42 0 0 5
1244 347
1244 337
1176 337
1176 663
1197 663
2 2 12 0 0 12416 0 35 39 0 0 5
1244 383
1244 400
1184 400
1184 523
1197 523
1 1 7 0 0 0 0 36 41 0 0 5
1196 346
1196 342
1181 342
1181 617
1197 617
1 0 13 0 0 4096 0 39 0 0 18 2
1197 514
1187 514
2 1 13 0 0 8320 0 36 40 0 0 4
1196 382
1187 382
1187 561
1197 561
2 0 5 0 0 0 0 41 0 0 20 2
1197 635
1141 635
1 4 5 0 0 0 0 37 39 0 0 6
1273 700
1306 700
1306 714
1141 714
1141 541
1197 541
2 0 14 0 0 4096 0 42 0 0 22 2
1197 681
1158 681
2 4 14 0 0 8320 0 37 40 0 0 4
1237 700
1158 700
1158 588
1197 588
3 0 15 0 0 8320 0 43 0 0 33 5
1305 635
1308 635
1308 538
1286 538
1286 488
4 0 16 0 0 12416 0 38 0 0 34 4
1304 574
1304 547
1275 547
1275 470
3 2 17 0 0 4224 0 42 43 0 0 3
1242 672
1242 644
1259 644
3 1 18 0 0 4224 0 41 43 0 0 2
1242 626
1259 626
5 2 19 0 0 4224 0 40 38 0 0 2
1242 574
1259 574
5 1 20 0 0 4224 0 39 38 0 0 3
1242 527
1242 565
1258 565
3 0 21 0 0 4096 0 46 0 0 36 2
1241 454
1301 454
3 2 22 0 0 4224 0 48 47 0 0 3
1350 525
1350 497
1367 497
3 1 23 0 0 4224 0 49 47 0 0 2
1350 479
1367 479
0 1 24 0 0 12416 0 0 48 35 0 5
1315 423
1315 438
1291 438
1291 516
1305 516
2 2 15 0 0 0 0 49 45 0 0 4
1305 488
1249 488
1249 432
1262 432
1 1 16 0 0 0 0 49 45 0 0 4
1305 470
1254 470
1254 414
1262 414
3 1 24 0 0 0 0 45 44 0 0 2
1311 423
1346 423
2 2 21 0 0 8320 0 48 44 0 0 4
1305 534
1301 534
1301 441
1346 441
1 3 25 0 0 4224 0 15 23 0 0 5
1553 270
1553 725
1124 725
1124 432
1097 432
1 0 26 0 0 8320 0 2 0 0 54 7
152 990
152 959
1021 959
1021 737
1026 737
1026 706
1008 706
1 3 27 0 0 8320 0 7 29 0 0 9
150 887
150 851
1034 851
1034 737
1039 737
1039 599
950 599
950 583
960 583
0 0 7 0 0 0 0 0 0 6 50 2
891 273
891 342
0 0 8 0 0 0 0 0 0 7 48 2
900 246
900 337
0 0 9 0 0 0 0 0 0 8 46 2
909 228
909 332
3 1 28 0 0 8320 0 52 21 0 0 9
817 488
845 488
845 290
1030 290
1030 393
966 393
966 407
898 407
898 445
2 2 29 0 0 12416 0 33 21 0 0 6
992 384
962 384
962 404
894 404
894 463
898 463
3 0 9 0 0 0 0 28 0 0 46 2
899 532
873 532
1 3 9 0 0 0 0 33 27 0 0 5
992 348
992 332
873 332
873 579
899 579
2 0 8 0 0 0 0 27 0 0 48 2
899 570
878 570
1 1 8 0 0 0 0 32 25 0 0 5
946 347
946 337
878 337
878 663
899 663
2 2 30 0 0 12416 0 32 28 0 0 5
946 383
946 400
886 400
886 523
899 523
1 1 7 0 0 0 0 31 26 0 0 5
898 346
898 342
883 342
883 617
899 617
1 0 31 0 0 4096 0 28 0 0 52 2
899 514
889 514
2 1 31 0 0 8320 0 31 27 0 0 4
898 382
889 382
889 561
899 561
2 0 26 0 0 0 0 26 0 0 54 2
899 635
836 635
1 4 26 0 0 0 0 30 28 0 0 6
975 700
1008 700
1008 714
836 714
836 541
899 541
2 0 32 0 0 4096 0 25 0 0 56 2
899 681
859 681
2 4 32 0 0 8320 0 30 27 0 0 4
939 700
859 700
859 588
899 588
3 0 33 0 0 8320 0 24 0 0 67 5
1007 635
1010 635
1010 538
988 538
988 488
4 0 34 0 0 12416 0 29 0 0 68 4
1006 574
1006 547
977 547
977 470
3 2 35 0 0 4224 0 25 24 0 0 3
944 672
944 644
961 644
3 1 36 0 0 4224 0 26 24 0 0 2
944 626
961 626
5 2 37 0 0 4224 0 27 29 0 0 2
944 574
961 574
5 1 38 0 0 4224 0 28 29 0 0 3
944 527
944 565
960 565
3 0 39 0 0 4096 0 21 0 0 70 2
943 454
1003 454
3 2 40 0 0 4224 0 19 20 0 0 3
1052 525
1052 497
1069 497
3 1 41 0 0 4224 0 18 20 0 0 2
1052 479
1069 479
0 1 42 0 0 12416 0 0 19 69 0 5
1017 423
1017 438
993 438
993 516
1007 516
2 2 33 0 0 0 0 18 22 0 0 4
1007 488
951 488
951 432
964 432
1 1 34 0 0 0 0 18 22 0 0 4
1007 470
956 470
956 414
964 414
3 1 42 0 0 0 0 22 23 0 0 2
1013 423
1048 423
2 2 39 0 0 8320 0 19 23 0 0 4
1007 534
1003 534
1003 441
1048 441
1 3 43 0 0 8320 0 14 55 0 0 5
1579 269
1579 734
826 734
826 432
799 432
1 0 44 0 0 8320 0 3 0 0 88 7
188 991
188 971
723 971
723 737
728 737
728 706
710 706
1 3 45 0 0 8320 0 6 61 0 0 9
186 888
186 858
736 858
736 737
741 737
741 599
652 599
652 583
662 583
0 0 7 0 0 0 0 0 0 6 84 2
593 273
593 342
0 0 8 0 0 0 0 0 0 7 82 2
602 246
602 337
0 0 9 0 0 0 0 0 0 8 80 2
611 228
611 332
3 1 46 0 0 8320 0 79 53 0 0 9
519 488
547 488
547 288
732 288
732 393
668 393
668 407
600 407
600 445
2 2 47 0 0 12416 0 65 53 0 0 6
694 384
664 384
664 404
596 404
596 463
600 463
3 0 9 0 0 0 0 60 0 0 80 2
601 532
575 532
1 3 9 0 0 0 0 65 59 0 0 5
694 348
694 332
575 332
575 579
601 579
2 0 8 0 0 0 0 59 0 0 82 2
601 570
580 570
1 1 8 0 0 0 0 64 57 0 0 5
648 347
648 337
580 337
580 663
601 663
2 2 48 0 0 12416 0 64 60 0 0 5
648 383
648 400
588 400
588 523
601 523
1 1 7 0 0 0 0 63 58 0 0 5
600 346
600 342
585 342
585 617
601 617
1 0 49 0 0 4096 0 60 0 0 86 2
601 514
591 514
2 1 49 0 0 8320 0 63 59 0 0 4
600 382
591 382
591 561
601 561
2 0 44 0 0 0 0 58 0 0 88 2
601 635
549 635
1 4 44 0 0 0 0 62 60 0 0 6
677 700
710 700
710 714
549 714
549 541
601 541
2 0 50 0 0 4096 0 57 0 0 90 2
601 681
566 681
2 4 50 0 0 8320 0 62 59 0 0 4
641 700
566 700
566 588
601 588
3 0 51 0 0 8320 0 56 0 0 101 5
709 635
712 635
712 538
690 538
690 488
4 0 52 0 0 12416 0 61 0 0 102 4
708 574
708 547
679 547
679 470
3 2 53 0 0 4224 0 57 56 0 0 3
646 672
646 644
663 644
3 1 54 0 0 4224 0 58 56 0 0 2
646 626
663 626
5 2 55 0 0 4224 0 59 61 0 0 2
646 574
663 574
5 1 56 0 0 4224 0 60 61 0 0 3
646 527
646 565
662 565
3 0 57 0 0 4096 0 53 0 0 104 2
645 454
705 454
3 2 58 0 0 4224 0 51 52 0 0 3
754 525
754 497
771 497
3 1 59 0 0 4224 0 50 52 0 0 2
754 479
771 479
0 1 60 0 0 12416 0 0 51 103 0 5
719 423
719 438
695 438
695 516
709 516
2 2 51 0 0 0 0 50 54 0 0 4
709 488
653 488
653 432
666 432
1 1 52 0 0 0 0 50 54 0 0 4
709 470
658 470
658 414
666 414
3 1 60 0 0 0 0 54 55 0 0 2
715 423
750 423
2 2 57 0 0 8320 0 51 55 0 0 4
709 534
705 534
705 441
750 441
1 3 61 0 0 8320 0 13 76 0 0 5
1603 269
1603 743
528 743
528 432
501 432
1 0 62 0 0 12432 0 4 0 0 121 7
220 991
220 984
425 984
425 737
430 737
430 706
412 706
0 0 7 0 0 0 0 0 0 6 117 2
295 273
295 342
0 0 8 0 0 0 0 0 0 7 115 2
304 246
304 337
0 0 9 0 0 0 0 0 0 8 113 2
313 228
313 332
1 1 63 0 0 4224 0 9 78 0 0 8
220 788
220 319
434 319
434 393
370 393
370 407
302 407
302 445
2 2 64 0 0 12416 0 66 78 0 0 6
396 384
366 384
366 404
298 404
298 463
302 463
3 0 9 0 0 0 0 71 0 0 113 2
303 532
270 532
1 3 9 0 0 0 0 66 72 0 0 5
396 348
396 332
270 332
270 579
303 579
2 0 8 0 0 0 0 72 0 0 115 2
303 570
282 570
1 1 8 0 0 0 0 67 74 0 0 5
350 347
350 337
282 337
282 663
303 663
2 2 65 0 0 12416 0 67 71 0 0 5
350 383
350 400
290 400
290 523
303 523
1 1 7 0 0 0 0 68 73 0 0 5
302 346
302 342
287 342
287 617
303 617
1 0 66 0 0 4096 0 71 0 0 119 2
303 514
293 514
2 1 66 0 0 8320 0 68 72 0 0 4
302 382
293 382
293 561
303 561
2 0 62 0 0 0 0 73 0 0 121 2
303 635
244 635
1 4 62 0 0 0 0 69 71 0 0 6
379 700
412 700
412 714
244 714
244 541
303 541
2 0 67 0 0 4096 0 74 0 0 123 2
303 681
265 681
2 4 67 0 0 8320 0 69 72 0 0 4
343 700
265 700
265 588
303 588
3 0 68 0 0 8320 0 75 0 0 134 5
411 635
414 635
414 538
392 538
392 488
4 0 69 0 0 12416 0 70 0 0 135 4
410 574
410 547
381 547
381 470
3 2 70 0 0 4224 0 74 75 0 0 3
348 672
348 644
365 644
3 1 71 0 0 4224 0 73 75 0 0 2
348 626
365 626
5 2 72 0 0 4224 0 72 70 0 0 2
348 574
365 574
5 1 73 0 0 4224 0 71 70 0 0 3
348 527
348 565
364 565
3 0 74 0 0 4096 0 78 0 0 137 2
347 454
407 454
3 2 75 0 0 4224 0 80 79 0 0 3
456 525
456 497
473 497
3 1 76 0 0 4224 0 81 79 0 0 2
456 479
473 479
0 1 77 0 0 12416 0 0 80 136 0 5
421 423
421 438
397 438
397 516
411 516
2 2 68 0 0 0 0 81 77 0 0 4
411 488
355 488
355 432
368 432
1 1 69 0 0 0 0 81 77 0 0 4
411 470
360 470
360 414
368 414
3 1 77 0 0 0 0 77 76 0 0 2
417 423
452 423
2 2 74 0 0 8320 0 80 76 0 0 4
411 534
407 534
407 441
452 441
24
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
169 1009 206 1033
179 1017 195 1033
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
202 1008 239 1032
212 1016 228 1032
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
135 1008 172 1032
145 1016 161 1032
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
101 1007 138 1031
111 1015 127 1031
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
200 905 237 929
210 913 226 929
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
168 906 205 930
178 914 194 930
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
133 905 170 929
143 913 159 929
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
99 904 136 928
109 912 125 928
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
983 575 1020 599
993 583 1009 599
2 X0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
988 636 1025 660
998 644 1014 660
2 Y0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
924 452 961 476
934 460 950 476
2 Z0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1222 452 1259 476
1232 460 1248 476
2 Z0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1286 636 1323 660
1296 644 1312 660
2 Y0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1281 575 1318 599
1291 583 1307 599
2 X0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
685 575 722 599
695 583 711 599
2 X0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
690 636 727 660
700 644 716 660
2 Y0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
626 452 663 476
636 460 652 476
2 Z0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
328 452 365 476
338 460 354 476
2 Z0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
392 636 429 660
402 644 418 660
2 Y0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
387 575 424 599
397 583 413 599
2 X0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
101 804 138 828
111 812 127 828
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
135 805 172 829
145 813 161 829
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
170 806 207 830
180 814 196 830
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
202 805 263 829
212 813 252 829
5 Count
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
