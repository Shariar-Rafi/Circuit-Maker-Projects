CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
540 0 30 100 10
216 93 1364 691
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
426 213 567 334
42991634 0
0
6 Title:
5 Name:
0
0
0
34
13 Logic Switch~
5 595 322 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44803.4 0
0
13 Logic Switch~
5 596 362 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44803.4 1
0
13 Logic Switch~
5 595 399 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44803.4 2
0
13 Logic Switch~
5 594 435 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
44803.4 3
0
13 Logic Switch~
5 595 698 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
44803.4 4
0
13 Logic Switch~
5 595 734 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
44803.4 5
0
13 Logic Switch~
5 592 771 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
44803.4 6
0
13 Logic Switch~
5 588 818 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
44803.4 7
0
13 Logic Switch~
5 725 283 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
44803.4 8
0
9 2-In XOR~
219 959 610 0 3 22
0 23 24 19
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
972 0 0
2
44803.4 9
0
9 2-In XOR~
219 1021 664 0 3 22
0 19 18 22
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1B
3 -26 24 -18
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3472 0 0
2
44803.4 10
0
9 2-In AND~
219 1112 720 0 3 22
0 19 18 21
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9998 0 0
2
44803.4 11
0
9 2-In AND~
219 1113 783 0 3 22
0 24 23 20
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3536 0 0
2
44803.4 12
0
14 Logic Display~
6 1533 285 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L23
-10 -22 11 -14
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
44803.4 13
0
8 2-In OR~
219 1206 719 0 3 22
0 21 20 5
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3835 0 0
2
44803.4 14
0
9 2-In XOR~
219 961 348 0 3 22
0 28 2 29
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3670 0 0
2
44803.4 15
0
9 2-In XOR~
219 1089 374 0 3 22
0 29 30 27
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U1D
3 -26 24 -18
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
5616 0 0
2
44803.4 16
0
9 2-In AND~
219 1114 458 0 3 22
0 30 29 26
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9323 0 0
2
44803.4 17
0
9 2-In AND~
219 1115 521 0 3 22
0 2 28 25
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
317 0 0
2
44803.4 18
0
14 Logic Display~
6 1572 289 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L21
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
44803.4 19
0
8 2-In OR~
219 1208 457 0 3 22
0 26 25 18
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
4299 0 0
2
44803.4 20
0
8 2-In OR~
219 1224 1066 0 3 22
0 15 14 4
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
9672 0 0
2
44803.4 21
0
14 Logic Display~
6 1483 285 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
44803.4 22
0
9 2-In AND~
219 1131 1130 0 3 22
0 3 17 14
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
6369 0 0
2
44803.4 23
0
9 2-In AND~
219 1130 1067 0 3 22
0 13 5 15
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9172 0 0
2
44803.4 24
0
9 2-In XOR~
219 1039 1011 0 3 22
0 13 5 16
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U5A
3 -26 24 -18
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7100 0 0
2
44803.4 25
0
9 2-In XOR~
219 977 957 0 3 22
0 17 3 13
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U5B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3820 0 0
2
44803.4 26
0
8 2-In OR~
219 1238 1456 0 3 22
0 9 8 7
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7678 0 0
2
44803.4 27
0
14 Logic Display~
6 1318 295 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
44803.4 28
0
14 Logic Display~
6 1441 289 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
44803.4 29
0
9 2-In AND~
219 1145 1520 0 3 22
0 12 11 8
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3409 0 0
2
44803.4 30
0
9 2-In AND~
219 1144 1457 0 3 22
0 6 4 9
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3951 0 0
2
44803.4 31
0
9 2-In XOR~
219 1053 1401 0 3 22
0 6 4 10
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U5C
3 -26 24 -18
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
8885 0 0
2
44803.4 32
0
9 2-In XOR~
219 991 1347 0 3 22
0 11 12 6
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U5D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3780 0 0
2
44803.4 33
0
45
1 2 2 0 0 8320 0 8 16 0 0 4
600 818
775 818
775 357
945 357
1 2 3 0 0 12416 0 6 27 0 0 4
607 734
619 734
619 966
961 966
3 2 4 0 0 8320 0 22 32 0 0 7
1257 1066
1257 1199
754 1199
754 1476
1112 1476
1112 1466
1120 1466
3 2 5 0 0 8320 0 15 25 0 0 9
1239 719
1239 832
745 832
745 949
746 949
746 1086
1098 1086
1098 1076
1106 1076
2 0 4 0 0 0 0 33 0 0 3 3
1037 1410
1022 1410
1022 1476
1 0 6 0 0 8192 0 33 0 0 7 3
1037 1392
1033 1392
1033 1347
3 1 6 0 0 8320 0 34 32 0 0 4
1024 1347
1099 1347
1099 1448
1120 1448
3 1 7 0 0 16512 0 28 29 0 0 6
1271 1456
1319 1456
1319 1473
1338 1473
1338 313
1318 313
3 2 8 0 0 8320 0 31 28 0 0 4
1166 1520
1217 1520
1217 1465
1225 1465
3 1 9 0 0 4224 0 32 28 0 0 4
1165 1457
1217 1457
1217 1447
1225 1447
3 1 10 0 0 16512 0 33 30 0 0 5
1086 1401
1247 1401
1247 1380
1441 1380
1441 307
0 2 11 0 0 4096 0 0 31 15 0 3
929 1334
929 1529
1121 1529
0 1 12 0 0 8192 0 0 31 14 0 3
961 1374
961 1511
1121 1511
1 2 12 0 0 8320 0 5 34 0 0 6
607 698
636 698
636 1374
967 1374
967 1356
975 1356
1 1 11 0 0 8320 0 1 34 0 0 6
607 322
708 322
708 1334
967 1334
967 1338
975 1338
2 0 5 0 0 0 0 26 0 0 4 3
1023 1020
1008 1020
1008 1086
1 0 13 0 0 8192 0 26 0 0 18 3
1023 1002
1019 1002
1019 957
3 1 13 0 0 8320 0 27 25 0 0 4
1010 957
1085 957
1085 1058
1106 1058
3 2 14 0 0 8320 0 24 22 0 0 4
1152 1130
1203 1130
1203 1075
1211 1075
3 1 15 0 0 4224 0 25 22 0 0 4
1151 1067
1203 1067
1203 1057
1211 1057
3 1 16 0 0 16512 0 26 23 0 0 5
1072 1011
1233 1011
1233 990
1483 990
1483 303
0 2 17 0 0 8192 0 0 24 24 0 3
908 944
908 1139
1107 1139
0 1 3 0 0 0 0 0 24 2 0 3
945 966
945 1121
1107 1121
1 1 17 0 0 8320 0 2 27 0 0 6
608 362
664 362
664 944
953 944
953 948
961 948
2 0 18 0 0 8192 0 11 0 0 28 3
1005 673
990 673
990 739
1 0 19 0 0 8192 0 11 0 0 27 3
1005 655
1001 655
1001 610
3 1 19 0 0 8320 0 10 12 0 0 4
992 610
1067 610
1067 711
1088 711
3 2 18 0 0 8320 0 21 12 0 0 7
1241 457
1241 556
746 556
746 739
1080 739
1080 729
1088 729
3 2 20 0 0 8320 0 13 15 0 0 4
1134 783
1185 783
1185 728
1193 728
3 1 21 0 0 4224 0 12 15 0 0 4
1133 720
1185 720
1185 710
1193 710
3 1 22 0 0 16512 0 11 14 0 0 5
1054 664
1215 664
1215 643
1533 643
1533 303
0 2 23 0 0 8192 0 0 13 35 0 3
878 597
878 792
1089 792
0 1 24 0 0 8320 0 0 13 34 0 3
894 637
894 774
1089 774
1 2 24 0 0 0 0 7 10 0 0 6
604 771
792 771
792 637
935 637
935 619
943 619
1 1 23 0 0 12416 0 3 10 0 0 6
607 399
633 399
633 597
935 597
935 601
943 601
3 2 25 0 0 8320 0 19 21 0 0 4
1136 521
1187 521
1187 466
1195 466
3 1 26 0 0 4224 0 18 21 0 0 4
1135 458
1187 458
1187 448
1195 448
3 1 27 0 0 12416 0 17 20 0 0 5
1122 374
1217 374
1217 381
1572 381
1572 307
0 2 28 0 0 8320 0 0 19 45 0 3
879 335
879 530
1091 530
0 1 2 0 0 0 0 0 19 1 0 5
906 357
906 375
905 375
905 512
1091 512
0 2 29 0 0 4224 0 0 18 44 0 3
1003 348
1003 467
1090 467
0 1 30 0 0 8192 0 0 18 43 0 3
1038 422
1038 449
1090 449
1 2 30 0 0 12416 0 9 17 0 0 6
737 283
828 283
828 422
1065 422
1065 383
1073 383
3 1 29 0 0 0 0 16 17 0 0 4
994 348
1065 348
1065 365
1073 365
1 1 28 0 0 0 0 4 16 0 0 7
606 435
606 488
731 488
731 335
937 335
937 339
945 339
82
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1178 726 1207 750
1188 734 1196 750
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1177 683 1206 707
1187 691 1195 707
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1234 698 1263 722
1244 706 1252 722
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1120 692 1149 716
1130 700 1138 716
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1075 723 1104 747
1085 731 1093 747
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1076 687 1105 711
1086 695 1094 711
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1121 757 1150 781
1131 765 1139 781
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1078 789 1107 813
1088 797 1096 813
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1076 752 1105 776
1086 760 1094 776
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1058 645 1087 669
1068 653 1076 669
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1057 596 1086 620
1067 604 1075 620
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1111 609 1140 633
1121 617 1129 633
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
975 580 1004 604
985 588 993 604
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
931 621 960 645
941 629 949 645
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
926 568 955 592
936 576 944 592
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1180 464 1209 488
1190 472 1198 488
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1179 421 1208 445
1189 429 1197 445
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1236 436 1265 460
1246 444 1254 460
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1122 430 1151 454
1132 438 1140 454
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1077 461 1106 485
1087 469 1095 485
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1078 425 1107 449
1088 433 1096 449
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1123 495 1152 519
1133 503 1141 519
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1080 527 1109 551
1090 535 1098 551
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1078 490 1107 514
1088 498 1096 514
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1060 383 1089 407
1070 391 1078 407
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1059 334 1088 358
1069 342 1077 358
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1113 347 1142 371
1123 355 1131 371
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
977 318 1006 342
987 326 995 342
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
933 359 962 383
943 367 951 383
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
928 306 957 330
938 314 946 330
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
944 915 973 939
954 923 962 939
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
949 968 978 992
959 976 967 992
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
993 927 1022 951
1003 935 1011 951
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1057 983 1086 1007
1067 991 1075 1007
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1019 968 1048 992
1029 976 1037 992
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1004 1030 1033 1054
1014 1038 1022 1054
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1094 1099 1123 1123
1104 1107 1112 1123
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1096 1136 1125 1160
1106 1144 1114 1160
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1139 1104 1168 1128
1149 1112 1157 1128
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1094 1034 1123 1058
1104 1042 1112 1058
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1093 1070 1122 1094
1103 1078 1111 1094
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1138 1039 1167 1063
1148 1047 1156 1063
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1252 1045 1281 1069
1262 1053 1270 1069
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1195 1030 1224 1054
1205 1038 1213 1054
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1196 1073 1225 1097
1206 1081 1214 1097
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1112 1264 1141 1288
1122 1272 1130 1288
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
958 1305 987 1329
968 1313 976 1329
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
963 1358 992 1382
973 1366 981 1382
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1007 1317 1036 1341
1017 1325 1025 1341
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1143 1346 1172 1370
1153 1354 1161 1370
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1089 1333 1118 1357
1099 1341 1107 1357
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1090 1382 1119 1406
1100 1390 1108 1406
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1108 1489 1137 1513
1118 1497 1126 1513
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1110 1526 1139 1550
1120 1534 1128 1550
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1153 1494 1182 1518
1163 1502 1171 1518
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1108 1424 1137 1448
1118 1432 1126 1448
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1107 1460 1136 1484
1117 1468 1125 1484
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1152 1429 1181 1453
1162 1437 1170 1453
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1266 1435 1295 1459
1276 1443 1284 1459
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1209 1420 1238 1444
1219 1428 1227 1444
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1210 1463 1239 1487
1220 1471 1228 1487
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
543 339 580 363
555 348 567 364
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
545 383 580 407
556 392 568 408
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
544 421 579 445
555 430 567 446
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
553 674 588 698
564 683 576 699
2 B4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
547 715 588 738
560 725 574 740
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
544 755 585 778
557 765 571 780
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
540 803 581 826
553 813 567 828
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
812 520 860 543
825 530 846 545
3 cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
813 801 859 824
825 811 846 826
3 cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
844 1168 890 1191
856 1178 877 1193
3 cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1288 248 1343 271
1301 258 1329 273
4 cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1412 236 1455 260
1419 240 1447 256
4 sum4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1456 233 1497 257
1462 238 1490 254
4 sum3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1507 233 1548 257
1513 238 1541 254
4 sum2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1546 238 1587 262
1552 242 1580 258
4 sum1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
542 310 571 334
549 314 563 330
2 A4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
654 273 697 297
661 278 689 294
4 C in
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 40
1008 111 1063 235
1014 116 1056 212
40 Cout=1

Sum1=0
Sum2=1
Sum3=1
Sum4=1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 42
769 97 847 181
776 101 839 165
42 A1=1 B1=1
A2=1 B2=1
A3=1 B3=1
A4=1 B4=1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
784 46 918 70
791 50 910 66
17 4 bit full adder:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
1382 37 1446 81
1389 41 1438 73
16 Group-5
_______
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
