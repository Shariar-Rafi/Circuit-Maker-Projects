CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
216 93 1364 691
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
426 213 567 334
42991634 0
0
6 Title:
5 Name:
0
0
0
19
6 74136~
219 302 477 0 3 22
0 3 2 7
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
5130 0 0
2
44803.5 18
0
6 74136~
219 305 424 0 3 22
0 4 2 8
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
391 0 0
2
44803.5 17
0
6 74136~
219 309 371 0 3 22
0 5 2 9
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U6C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
3124 0 0
2
44803.5 16
0
6 74136~
219 300 317 0 3 22
0 6 2 10
0
0 0 608 0
7 74LS136
-24 -24 25 -16
3 U6D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
3421 0 0
2
44803.5 15
0
14 Logic Display~
6 812 170 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
44803.5 14
0
14 Logic Display~
6 773 172 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
44803.5 13
0
14 Logic Display~
6 726 176 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
44803.5 12
0
14 Logic Display~
6 682 178 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
44803.5 11
0
14 Logic Display~
6 639 176 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
44803.5 10
0
6 74LS83
105 509 240 0 14 29
0 19 18 17 16 10 9 8 7 2
14 13 12 11 15
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U8
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
972 0 0
2
44803.5 9
0
13 Logic Switch~
5 244 552 0 1 11
0 2
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V32
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
44803.5 8
0
13 Logic Switch~
5 156 423 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V31
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
44803.5 7
0
13 Logic Switch~
5 157 477 0 1 11
0 3
0
0 0 21344 0
2 0V
-5 -16 9 -8
3 V30
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3536 0 0
2
44803.5 6
0
13 Logic Switch~
5 163 367 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V29
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4597 0 0
2
44803.5 5
0
13 Logic Switch~
5 164 331 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V28
-11 -27 10 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
44803.5 4
0
13 Logic Switch~
5 159 229 0 1 11
0 16
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V27
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3670 0 0
2
44803.5 3
0
13 Logic Switch~
5 159 190 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V26
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5616 0 0
2
44803.5 2
0
13 Logic Switch~
5 164 153 0 1 11
0 18
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V25
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9323 0 0
2
44803.5 1
0
13 Logic Switch~
5 163 120 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V24
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
317 0 0
2
44803.5 0
0
22
0 9 2 0 0 16 0 0 10 9 0 4
265 526
449 526
449 285
477 285
0 2 2 0 0 16 0 0 1 9 0 2
265 486
286 486
1 1 3 0 0 16 0 13 1 0 0 4
169 477
278 477
278 468
286 468
0 2 2 0 0 16 0 0 2 9 0 2
265 433
289 433
1 1 4 0 0 16 0 12 2 0 0 4
168 423
281 423
281 415
289 415
0 2 2 0 0 16 0 0 3 9 0 2
265 380
293 380
1 1 5 0 0 16 0 14 3 0 0 4
175 367
285 367
285 362
293 362
1 1 6 0 0 16 0 15 4 0 0 5
176 331
176 311
276 311
276 308
284 308
2 1 2 0 0 16 0 4 11 0 0 4
284 326
265 326
265 552
256 552
3 8 7 0 0 16 0 1 10 0 0 4
335 477
469 477
469 267
477 267
3 7 8 0 0 16 0 2 10 0 0 4
338 424
464 424
464 258
477 258
3 6 9 0 0 16 0 3 10 0 0 4
342 371
459 371
459 249
477 249
3 5 10 0 0 16 0 4 10 0 0 6
333 317
334 317
334 331
454 331
454 240
477 240
13 1 11 0 0 16 0 10 5 0 0 3
541 258
812 258
812 188
12 1 12 0 0 16 0 10 6 0 0 3
541 249
773 249
773 190
11 1 13 0 0 16 0 10 7 0 0 3
541 240
726 240
726 194
10 1 14 0 0 16 0 10 8 0 0 3
541 231
682 231
682 196
14 1 15 0 0 16 0 10 9 0 0 3
541 285
639 285
639 194
1 4 16 0 0 16 0 16 10 0 0 4
171 229
469 229
469 231
477 231
1 3 17 0 0 16 0 17 10 0 0 4
171 190
459 190
459 222
477 222
1 2 18 0 0 16 0 18 10 0 0 4
176 153
464 153
464 213
477 213
1 1 19 0 0 16 0 19 10 0 0 4
175 120
469 120
469 204
477 204
27
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
183 528 219 552
190 533 211 549
3 cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
435 17 548 59
443 22 539 52
27 4 bit adder 
substractor:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
842 362 951 386
852 370 940 386
11 which is 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
691 364 856 388
701 372 845 388
18 Subtarctor: 10-8=2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
98 410 135 434
108 418 124 434
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
106 210 143 234
116 218 132 234
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
105 315 142 339
115 323 131 339
2 B4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
104 363 141 387
114 371 130 387
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
102 460 139 484
112 468 128 484
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
105 106 142 130
115 114 131 130
2 A4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
105 140 142 164
115 148 131 164
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
105 176 142 200
115 184 131 200
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
328 301 365 325
338 309 354 325
2 11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
262 283 299 307
272 291 288 307
2 12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
262 320 299 344
272 328 288 344
2 13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
329 345 358 369
339 353 347 369
1 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
278 336 307 360
288 344 296 360
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
277 376 306 400
287 384 295 400
1 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
326 398 355 422
336 406 344 422
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
263 394 292 418
273 402 281 418
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
272 426 301 450
282 434 290 450
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
322 452 351 476
332 460 340 476
1 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
266 443 295 467
276 451 284 467
1 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
270 481 299 505
280 489 288 505
1 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
688 314 837 338
698 322 826 338
16 Adder: 10+10 =20
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
828 312 961 336
838 320 950 336
14 which is 10100
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
1662 1550 1735 1592
1670 1555 1726 1585
16 Group-5
_______
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
