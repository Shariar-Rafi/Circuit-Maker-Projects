CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 130 30 120 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
77 E:\Software (Installed and Running)\Electronics\CircuitMaker 2000 SP1\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
16
14 Logic Display~
6 468 156 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5130 0 0
2
44859.4 0
0
14 Logic Display~
6 440 157 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
391 0 0
2
44859.4 0
0
14 Logic Display~
6 414 157 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3124 0 0
2
44859.4 0
0
14 Logic Display~
6 382 157 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3421 0 0
2
44859.4 0
0
13 Logic Switch~
5 71 693 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8157 0 0
2
44859.4 0
0
14 Logic Display~
6 321 156 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
44859.4 0
0
13 Logic Switch~
5 18 433 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8901 0 0
2
44859.4 0
0
13 Logic Switch~
5 20 401 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7361 0 0
2
44859.4 0
0
13 Logic Switch~
5 20 369 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4747 0 0
2
44859.4 0
0
13 Logic Switch~
5 20 338 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
972 0 0
2
44859.4 0
0
13 Logic Switch~
5 20 308 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3472 0 0
2
44859.4 0
0
13 Logic Switch~
5 20 281 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9998 0 0
2
44859.4 0
0
13 Logic Switch~
5 20 252 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3536 0 0
2
44859.4 0
0
13 Logic Switch~
5 21 221 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4597 0 0
2
44859.4 0
0
13 Logic Switch~
5 19 188 0 1 11
0 0
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3835 0 0
2
44859.4 0
0
6 74LS83
105 278 284 0 1 29
0 0
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 0 0 0 0
1 U
3670 0 0
2
44859.4 0
0
14
13 1 0 0 0 0 0 16 1 0 0 3
310 302
468 302
468 174
12 1 0 0 0 0 0 16 2 0 0 3
310 293
440 293
440 175
11 1 0 0 0 0 0 16 3 0 0 3
310 284
414 284
414 175
10 1 0 0 0 0 0 16 4 0 0 3
310 275
382 275
382 175
14 1 0 0 0 0 0 16 6 0 0 3
310 329
321 329
321 174
1 9 0 0 0 0 0 7 16 0 0 4
30 433
248 433
248 329
246 329
1 8 0 0 0 0 0 8 16 0 0 4
32 401
242 401
242 311
246 311
1 7 0 0 0 0 0 9 16 0 0 4
32 369
236 369
236 302
246 302
1 6 0 0 0 0 0 10 16 0 0 5
32 338
32 324
233 324
233 293
246 293
1 5 0 0 0 16 0 11 16 0 0 5
32 308
32 288
238 288
238 284
246 284
1 4 0 0 0 0 0 12 16 0 0 5
32 281
32 274
238 274
238 275
246 275
1 3 0 0 0 0 0 13 16 0 0 5
32 252
32 262
238 262
238 266
246 266
1 2 0 0 0 0 0 14 16 0 0 4
33 221
233 221
233 257
246 257
1 1 0 0 0 0 0 15 16 0 0 4
31 188
238 188
238 248
246 248
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
