CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
216 93 1364 691
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
426 213 567 334
42991634 0
0
6 Title:
5 Name:
0
0
0
43
13 Logic Switch~
5 296 231 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6866 0 0
2
44817.4 1
0
13 Logic Switch~
5 296 281 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7670 0 0
2
44817.4 0
0
13 Logic Switch~
5 124 1869 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
951 0 0
2
44817.4 0
0
13 Logic Switch~
5 998 1678 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9536 0 0
2
44817.4 1
0
13 Logic Switch~
5 710 1689 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5495 0 0
2
44817.4 2
0
13 Logic Switch~
5 421 1702 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8152 0 0
2
44817.4 3
0
13 Logic Switch~
5 132 1714 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6223 0 0
2
44817.4 4
0
5 4030~
219 832 200 0 3 22
0 8 7 4
0
0 0 624 90
4 4030
-7 -24 21 -16
3 U5A
26 -3 47 5
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
5441 0 0
2
44817.4 12
0
5 4030~
219 643 190 0 3 22
0 8 9 5
0
0 0 624 90
4 4030
-7 -24 21 -16
3 U5B
26 -3 47 5
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
3189 0 0
2
44817.4 11
0
5 4030~
219 477 205 0 3 22
0 8 10 6
0
0 0 624 90
4 4030
-7 -24 21 -16
3 U5C
26 -3 47 5
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
8460 0 0
2
44817.4 10
0
7 Pulser~
4 248 355 0 10 12
0 30 31 11 32 0 0 10 10 1
8
0
0 0 4656 0
0
2 V6
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5179 0 0
2
44817.4 9
0
14 Logic Display~
6 836 118 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3593 0 0
2
44817.4 8
0
14 Logic Display~
6 646 126 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3928 0 0
2
44817.4 7
0
14 Logic Display~
6 482 134 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
363 0 0
2
44817.4 6
0
6 74112~
219 790 385 0 7 32
0 3 3 9 3 3 2 7
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U6A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 6 0
1 U
8132 0 0
2
44817.4 5
0
6 74112~
219 621 391 0 7 32
0 3 3 10 3 3 33 9
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U6B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 6 0
1 U
65 0 0
2
44817.4 4
0
6 74112~
219 441 394 0 7 32
0 3 3 11 3 3 34 10
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U7A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 7 0
1 U
6609 0 0
2
44817.4 3
0
12 Hex Display~
7 952 101 0 16 19
10 6 5 4 35 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
8995 0 0
2
44817.4 2
0
5 4023~
219 471 2074 0 4 22
0 14 13 16 17
0
0 0 624 0
4 4023
-14 -28 14 -20
4 U12B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 2 11 0
1 U
3918 0 0
2
44817.4 7
0
9 Inverter~
13 400 2091 0 2 22
0 21 13
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
7519 0 0
2
44817.4 8
0
9 Inverter~
13 406 2052 0 2 22
0 19 14
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
377 0 0
2
44817.4 9
0
9 Inverter~
13 408 1998 0 2 22
0 16 15
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
8816 0 0
2
44817.4 10
0
5 4023~
219 513 1972 0 4 22
0 21 19 15 18
0
0 0 624 0
4 4023
-14 -28 14 -20
4 U12A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 11 0
1 U
3877 0 0
2
44817.4 11
0
5 SCOPE
12 1164 1714 0 1 11
0 19
0
0 0 57584 0
3 TP8
-11 -4 10 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
926 0 0
2
44817.4 12
0
5 SCOPE
12 873 1726 0 1 11
0 20
0
0 0 57584 0
3 TP7
-11 -4 10 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7262 0 0
2
44817.4 13
0
5 SCOPE
12 594 1738 0 1 11
0 21
0
0 0 57584 0
3 TP6
-11 -4 10 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5267 0 0
2
44817.4 14
0
5 SCOPE
12 306 1749 0 1 11
0 22
0
0 0 57584 0
3 TP5
-11 -4 10 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8838 0 0
2
44817.4 15
0
5 SCOPE
12 145 1792 0 1 11
0 12
0
0 0 57584 0
3 TP4
-11 -4 10 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7159 0 0
2
44817.4 16
0
12 Hex Display~
7 1264 1741 0 18 19
10 22 21 20 19 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5812 0 0
2
44817.4 17
0
9 2-In XOR~
219 983 1750 0 3 22
0 20 16 25
0
0 0 624 0
5 74F86
-18 -24 17 -16
4 U11C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
331 0 0
2
44817.4 18
0
9 2-In XOR~
219 673 1763 0 3 22
0 21 16 24
0
0 0 624 0
5 74F86
-18 -24 17 -16
4 U11B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
9604 0 0
2
44817.4 19
0
9 2-In XOR~
219 380 1767 0 3 22
0 22 16 23
0
0 0 624 0
5 74F86
-18 -24 17 -16
4 U11A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
7518 0 0
2
44817.4 20
0
14 Logic Display~
6 1183 1591 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4832 0 0
2
44817.4 21
0
6 74112~
219 1111 1761 0 7 32
0 17 26 25 26 18 36 19
0
0 0 4720 0
5 74112
4 -60 39 -52
4 U10A
19 -61 47 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 9 0
1 U
6798 0 0
2
44817.4 22
0
14 Logic Display~
6 895 1593 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3336 0 0
2
44817.4 23
0
6 74112~
219 823 1772 0 7 32
0 17 27 24 27 18 37 20
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U8B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 8 0
1 U
8370 0 0
2
44817.4 24
0
6 74112~
219 534 1785 0 7 32
0 17 28 23 28 18 38 21
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U8A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 8 0
1 U
3910 0 0
2
44817.4 25
0
14 Logic Display~
6 616 1594 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
316 0 0
2
44817.4 26
0
14 Logic Display~
6 326 1593 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
536 0 0
2
44817.4 27
0
7 Pulser~
4 41 1811 0 10 12
0 12 39 12 40 0 0 10 10 1
8
0
0 0 4656 0
0
3 V13
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4460 0 0
2
44817.4 28
0
6 74112~
219 245 1797 0 7 32
0 17 29 12 29 18 41 22
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U7B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 7 0
1 U
3260 0 0
2
44817.4 29
0
5 SCOPE
12 665 1948 0 1 11
0 18
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5156 0 0
2
44817.4 30
0
5 SCOPE
12 665 2062 0 1 11
0 17
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3133 0 0
2
44817.4 31
0
80
6 0 2 0 0 4224 0 15 0 0 0 2
820 367
820 368
0 0 3 0 0 4096 0 0 0 0 16 2
613 400
613 403
0 3 4 0 0 4224 0 0 18 10 0 3
835 142
949 142
949 125
0 2 5 0 0 4224 0 0 18 12 0 3
646 152
955 152
955 125
0 1 6 0 0 4224 0 0 18 13 0 3
480 160
961 160
961 125
7 2 7 0 0 8320 0 15 8 0 0 3
814 349
844 349
844 219
0 1 8 0 0 4224 0 0 8 8 0 3
637 229
826 229
826 219
1 0 8 0 0 0 0 9 0 0 9 3
637 209
637 231
470 231
1 1 8 0 0 0 0 1 10 0 0 3
308 231
471 231
471 224
1 3 4 0 0 0 0 12 8 0 0 3
836 136
835 136
835 170
2 0 9 0 0 4224 0 9 0 0 18 2
655 209
655 358
3 1 5 0 0 0 0 9 13 0 0 4
646 160
646 162
646 162
646 144
3 1 6 0 0 0 0 10 14 0 0 3
480 175
480 152
482 152
2 7 10 0 0 12288 0 10 17 0 0 5
489 224
489 269
496 269
496 358
465 358
0 1 3 0 0 4096 0 0 15 25 0 3
766 298
790 298
790 322
0 5 3 0 0 8192 0 0 16 27 0 4
597 309
551 309
551 403
621 403
0 1 3 0 0 0 0 0 16 27 0 3
597 302
621 302
621 328
7 3 9 0 0 0 0 16 15 0 0 3
645 355
645 358
760 358
0 3 10 0 0 4224 0 0 16 14 0 4
496 356
586 356
586 364
591 364
3 3 11 0 0 12416 0 11 17 0 0 4
272 346
331 346
331 367
411 367
0 5 3 0 0 8192 0 0 15 25 0 5
766 290
731 290
731 407
790 407
790 397
0 5 3 0 0 0 0 0 17 23 0 4
441 299
357 299
357 406
441 406
0 1 3 0 0 0 0 0 17 27 0 3
442 281
441 281
441 331
0 4 3 0 0 0 0 0 15 25 0 4
766 309
746 309
746 367
766 367
0 2 3 0 0 4096 0 0 15 27 0 3
596 281
766 281
766 349
0 4 3 0 0 0 0 0 16 27 0 4
597 319
568 319
568 373
597 373
0 2 3 0 0 4224 0 0 16 29 0 3
417 281
597 281
597 355
0 4 3 0 0 0 0 0 17 29 0 4
417 329
385 329
385 376
417 376
1 2 3 0 0 0 0 2 17 0 0 3
308 281
417 281
417 358
1 0 12 0 0 4096 0 28 0 0 32 2
145 1804
145 1802
1 0 12 0 0 12288 0 40 0 0 32 5
17 1802
7 1802
7 1788
103 1788
103 1802
3 3 12 0 0 4224 0 40 41 0 0 4
65 1802
207 1802
207 1770
215 1770
2 2 13 0 0 8320 0 20 19 0 0 3
421 2091
421 2074
447 2074
2 1 14 0 0 12416 0 21 19 0 0 4
427 2052
425 2052
425 2065
447 2065
2 3 15 0 0 4224 0 22 23 0 0 4
429 1998
487 1998
487 1981
489 1981
0 1 16 0 0 8192 0 0 22 62 0 3
247 1869
247 1998
393 1998
1 0 17 0 0 0 0 43 0 0 52 2
665 2074
665 2074
1 0 18 0 0 4096 0 42 0 0 57 4
665 1960
665 1987
664 1987
664 1985
1 0 19 0 0 4096 0 24 0 0 69 2
1164 1726
1164 1725
1 0 20 0 0 4096 0 25 0 0 72 2
873 1738
873 1736
1 0 21 0 0 4096 0 26 0 0 75 2
594 1750
594 1749
1 0 22 0 0 0 0 27 0 0 78 2
306 1761
306 1761
0 1 19 0 0 8192 0 0 21 58 0 5
308 1972
308 2036
374 2036
374 2052
391 2052
0 1 21 0 0 8192 0 0 20 59 0 4
382 1925
321 1925
321 2091
385 2091
0 1 22 0 0 4224 0 0 29 78 0 4
325 1634
1320 1634
1320 1765
1273 1765
0 2 21 0 0 4224 0 0 29 75 0 5
616 1642
1296 1642
1296 1783
1267 1783
1267 1765
0 3 20 0 0 8320 0 0 29 72 0 6
895 1627
895 1623
1288 1623
1288 1798
1261 1798
1261 1765
4 0 19 0 0 16384 0 29 0 0 69 6
1255 1765
1245 1765
1245 1822
1308 1822
1308 1610
1183 1610
0 1 17 0 0 4096 0 0 41 50 0 3
534 1649
245 1649
245 1734
0 1 17 0 0 0 0 0 37 51 0 3
823 1649
534 1649
534 1722
0 1 17 0 0 0 0 0 36 52 0 4
1111 1648
1111 1649
823 1649
823 1709
4 1 17 0 0 4224 0 19 34 0 0 5
498 2074
1233 2074
1233 1648
1111 1648
1111 1698
0 3 16 0 0 8192 0 0 19 62 0 4
193 1869
193 2109
447 2109
447 2083
0 5 18 0 0 4096 0 0 41 55 0 3
549 1810
245 1810
245 1809
0 5 18 0 0 0 0 0 37 56 0 4
824 1809
824 1810
534 1810
534 1797
0 5 18 0 0 0 0 0 36 57 0 3
1111 1809
823 1809
823 1784
4 5 18 0 0 8320 0 23 34 0 0 4
540 1972
540 1985
1111 1985
1111 1773
2 0 19 0 0 12416 0 23 0 0 69 5
489 1972
278 1972
278 1882
1179 1882
1179 1725
1 0 21 0 0 0 0 23 0 0 75 5
489 1963
382 1963
382 1893
583 1893
583 1749
0 2 16 0 0 4224 0 0 30 61 0 4
639 1869
962 1869
962 1759
967 1759
0 2 16 0 0 0 0 0 31 62 0 4
342 1869
641 1869
641 1772
657 1772
1 2 16 0 0 0 0 3 32 0 0 4
136 1869
344 1869
344 1776
364 1776
3 3 23 0 0 12416 0 32 37 0 0 4
413 1767
454 1767
454 1758
504 1758
3 3 24 0 0 4224 0 31 36 0 0 4
706 1763
788 1763
788 1745
793 1745
3 3 25 0 0 4224 0 30 34 0 0 3
1016 1750
1081 1750
1081 1734
1 1 20 0 0 0 0 35 30 0 0 4
895 1611
951 1611
951 1741
967 1741
1 1 21 0 0 0 0 38 31 0 0 3
616 1612
657 1612
657 1754
1 1 22 0 0 0 0 39 32 0 0 3
326 1611
364 1611
364 1758
1 7 19 0 0 0 0 33 34 0 0 3
1183 1609
1183 1725
1135 1725
0 4 26 0 0 4224 0 0 34 71 0 3
1050 1678
1050 1743
1087 1743
1 2 26 0 0 0 0 4 34 0 0 4
1010 1678
1072 1678
1072 1725
1087 1725
1 7 20 0 0 0 0 35 36 0 0 3
895 1611
895 1736
847 1736
0 4 27 0 0 4224 0 0 36 74 0 3
762 1689
762 1754
799 1754
1 2 27 0 0 0 0 5 36 0 0 4
722 1689
784 1689
784 1736
799 1736
1 7 21 0 0 0 0 38 37 0 0 3
616 1612
616 1749
558 1749
0 4 28 0 0 4224 0 0 37 77 0 3
473 1702
473 1767
510 1767
1 2 28 0 0 0 0 6 37 0 0 4
433 1702
495 1702
495 1749
510 1749
1 7 22 0 0 0 0 39 41 0 0 5
326 1611
326 1634
325 1634
325 1761
269 1761
0 4 29 0 0 4224 0 0 41 80 0 3
184 1714
184 1779
221 1779
1 2 29 0 0 0 0 7 41 0 0 4
144 1714
206 1714
206 1761
221 1761
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
259 267 290 290
266 272 282 287
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
264 211 287 234
271 216 279 231
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
191 163 256 243
199 168 247 228
25 S=1
(Down)
S=0 
(Up)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
160 26 279 68
167 31 271 61
25 Mod 8 up-down 
counter:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
1137 7 1210 49
1145 12 1201 42
16 Group-5
_______
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
267 1551 315 1574
280 1561 301 1576
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1186 1548 1234 1571
1199 1558 1220 1573
3 MSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
458 1500 613 1524
469 1509 601 1525
22 MOD 10 Asynchronous Up
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
631 1501 696 1525
642 1510 684 1526
7 Counter
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
