CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 390 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 108 756 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V28
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90047e-315 0
0
13 Logic Switch~
5 204 614 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90047e-315 5.43969e-315
0
5 7474~
219 371 678 0 6 22
0 7 7 8 2 9 6
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U5A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
3124 0 0
2
5.90047e-315 5.49797e-315
0
5 7474~
219 511 660 0 6 22
0 7 6 8 2 10 5
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U5B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
3421 0 0
2
5.90047e-315 5.49926e-315
0
5 7474~
219 629 662 0 6 22
0 7 5 8 2 11 4
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U6A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
8157 0 0
2
5.90047e-315 5.50056e-315
0
5 7474~
219 724 656 0 6 22
0 7 4 8 2 12 3
0
0 0 4720 0
4 7474
7 -60 35 -52
3 U6B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 2 0
1 U
5572 0 0
2
5.90047e-315 5.50185e-315
0
7 Pulser~
4 204 708 0 10 12
0 8 2 8 13 0 0 5 5 1
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8901 0 0
2
5.90047e-315 5.50315e-315
0
14 Logic Display~
6 436 545 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
5.90047e-315 5.50444e-315
0
14 Logic Display~
6 574 542 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.90047e-315 5.50574e-315
0
14 Logic Display~
6 681 541 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.90047e-315 5.50703e-315
0
14 Logic Display~
6 804 543 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.90047e-315 5.50833e-315
0
23
2 0 2 0 0 8208 0 7 0 0 4 4
174 708
144 708
144 747
174 747
0 4 2 0 0 4096 0 0 5 3 0 4
630 724
630 682
629 682
629 674
0 4 2 0 0 4224 0 0 6 13 0 3
506 724
724 724
724 668
1 4 2 0 0 0 0 1 3 0 0 7
120 756
174 756
174 747
201 747
201 756
371 756
371 690
6 1 3 0 0 8320 0 6 11 0 0 3
748 620
804 620
804 561
0 1 4 0 0 4224 0 0 10 20 0 2
681 626
681 559
0 1 5 0 0 4224 0 0 9 21 0 2
574 624
574 560
0 1 6 0 0 4096 0 0 8 22 0 2
436 642
436 563
0 1 7 0 0 4096 0 0 5 12 0 2
629 585
629 599
0 1 7 0 0 0 0 0 4 12 0 2
511 585
511 597
0 1 7 0 0 4096 0 0 3 12 0 2
371 585
371 615
0 1 7 0 0 8320 0 0 6 23 0 4
306 614
306 585
724 585
724 593
0 4 2 0 0 0 0 0 4 4 0 5
371 736
506 736
506 685
511 685
511 672
0 4 2 0 0 0 0 0 3 0 0 3
370 685
370 690
371 690
1 0 8 0 0 12288 0 7 0 0 19 5
180 699
170 699
170 685
255 685
255 699
0 3 8 0 0 0 0 0 3 19 0 3
324 699
324 660
347 660
0 3 8 0 0 0 0 0 4 19 0 3
476 699
476 642
487 642
0 3 8 0 0 0 0 0 5 19 0 3
591 699
591 644
605 644
3 3 8 0 0 4224 0 7 6 0 0 4
228 699
692 699
692 638
700 638
6 2 4 0 0 0 0 5 6 0 0 4
653 626
692 626
692 620
700 620
6 2 5 0 0 0 0 4 5 0 0 4
535 624
597 624
597 626
605 626
6 2 6 0 0 4224 0 3 4 0 0 4
395 642
479 642
479 624
487 624
1 2 7 0 0 0 0 2 3 0 0 4
216 614
339 614
339 642
347 642
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
326 429 371 453
332 433 364 449
4 Sipo
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
